module layer5_1#(
    parameter DATA_WIDTH = 32,
    parameter WIDTH = 28
)(
  input  [DATA_WIDTH*16-1:0] i_data,
  input              clk, rst, valid_in,
  output [DATA_WIDTH*32-1:0] o_data,
  output             valid_out
);
  wire [DATA_WIDTH*16-1:0] i_CORE_IP1 [31:0];
  wire padding_valid, valid_in_pipeline2D, valid_in_bias;
  wire [31:0] counter_col, counter_row;
  wire [3:0] valid_pipeline2D;
  wire [4:0] valid_pipeline_bias;

/// CON2D_1///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011011011000001111001000),
      .k2(32'b00111101101000110011101100010100),
      .k3(32'b00111101001111111111011111010010),
      .k4(32'b00111101101000011101011000011001),
      .k5(32'b10111101101101101001011000000100),
      .k6(32'b00111101000100111111100011001100),
      .k7(32'b10111101001100111000000000010011),
      .k8(32'b00111101001010111001110011011001),
      .k9(32'b00111100001101101101011101110101)
  ) CON2D_1(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100000100110101001000111),
      .k2(32'b00111101001101111101000001010110),
      .k3(32'b00111100111111011000101000000111),
      .k4(32'b00111101111100101011001011101010),
      .k5(32'b00111101100010010001100010001011),
      .k6(32'b10111101000011011011111101001101),
      .k7(32'b00111101110001000100101011001011),
      .k8(32'b00111101101010011101001101010010),
      .k9(32'b10111101100100000001010001001000)
  ) CON2D_2(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111110110100100010010000),
      .k2(32'b10111101001000001011101111111111),
      .k3(32'b10111101110100000001000100011000),
      .k4(32'b00111101000101000000001110110101),
      .k5(32'b10111101001110100111000000000010),
      .k6(32'b10111101100010001001111101000100),
      .k7(32'b10111101110001110010000110011000),
      .k8(32'b00111101111110001100011100010101),
      .k9(32'b10111101011110000011000100101100)
  ) CON2D_3(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111000001001010111100),
      .k2(32'b00111101100100011001010101000000),
      .k3(32'b00111010011001001100111111100100),
      .k4(32'b00111101110011011010001000111110),
      .k5(32'b00111010111111101000101101100100),
      .k6(32'b10111101100000111110011111100101),
      .k7(32'b10111101100101101111111011111011),
      .k8(32'b10111101101000011000101000010010),
      .k9(32'b00111101000100010010010000100000)
  ) CON2D_4(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100001100111100001111001),
      .k2(32'b00111101110001010101001010010100),
      .k3(32'b10111101101000010110110111010011),
      .k4(32'b00111101111100001010110100111111),
      .k5(32'b10111101100101100010010010111011),
      .k6(32'b00111101110011100110011101000111),
      .k7(32'b10111100011100011011001111011011),
      .k8(32'b00111101101000001000001011010001),
      .k9(32'b00111101101110101111111110001001)
  ) CON2D_5(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100001101111011011001011111),
      .k2(32'b10111101000110100111100010001111),
      .k3(32'b00111101010000001011010100011101),
      .k4(32'b00111101101111001011001111110100),
      .k5(32'b00111100001110001110110100011111),
      .k6(32'b10111101111100001110010101111111),
      .k7(32'b00111100010101010101101000000011),
      .k8(32'b10111100100011100101000011111101),
      .k9(32'b00111101011001000101101100001111)
  ) CON2D_6(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011101110101100100000100110),
      .k2(32'b00111010111001010111000111001101),
      .k3(32'b00111101100000111010111101100011),
      .k4(32'b10111101010011001111011001110110),
      .k5(32'b00111101111111000010101101110010),
      .k6(32'b00111101110100000111010011001101),
      .k7(32'b00111101100000011110001100001001),
      .k8(32'b10111011101010101011100101000000),
      .k9(32'b00111010110101111100111010110010)
  ) CON2D_7(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111110111111100011101),
      .k2(32'b00111001110001000011111111111101),
      .k3(32'b00111100110100010000111000001000),
      .k4(32'b00111101111000101000111010011010),
      .k5(32'b10111101111000011111000110110000),
      .k6(32'b10111100101000000111010101011111),
      .k7(32'b10111100101111110111010001000100),
      .k8(32'b10111101110001000111100000100101),
      .k9(32'b00111100000100001101110110011100)
  ) CON2D_8(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000000100011001011110010),
      .k2(32'b00111101001111000011000111101010),
      .k3(32'b10111101000001001000010010110010),
      .k4(32'b00111100100001100011000001001001),
      .k5(32'b10111101101011001011010101011100),
      .k6(32'b10111101000000101000111000101000),
      .k7(32'b00111101001010111000010000011111),
      .k8(32'b00111101110010110110101100100000),
      .k9(32'b10111101110111000000010111110010)
  ) CON2D_9(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101001100000100111011101),
      .k2(32'b10111010101100101101111010100101),
      .k3(32'b00111100001100001001001000100110),
      .k4(32'b10111101100101111100010011101000),
      .k5(32'b00111100101101101101111111111001),
      .k6(32'b10111100110000111100010110000011),
      .k7(32'b00111101001110011111001010101101),
      .k8(32'b00111100000101001011011101010110),
      .k9(32'b00111100100010001100010101011001)
  ) CON2D_10(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111000010001100001010100),
      .k2(32'b10111100001001110111101101100111),
      .k3(32'b10111011010111110010000100001011),
      .k4(32'b10111101101100110101101101110100),
      .k5(32'b10111100001000001011100101001110),
      .k6(32'b10111101111101100110001111001111),
      .k7(32'b00111011110011001101111100111101),
      .k8(32'b00111101001001100111111001011000),
      .k9(32'b00111011101000000000100111101111)
  ) CON2D_11(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111000101110101011010110101000),
      .k2(32'b00111101101011100011001000101110),
      .k3(32'b10111101110101101101101010110101),
      .k4(32'b00111101000100010110001000101010),
      .k5(32'b10111100111100100010001001100000),
      .k6(32'b10111101101000000011001111000100),
      .k7(32'b10111101101011100110001011100000),
      .k8(32'b10111101011011100101110011111100),
      .k9(32'b00111100011101010011100111011101)
  ) CON2D_12(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100100011111010000001110),
      .k2(32'b10111101100000010000100100110011),
      .k3(32'b00111101100101010111010101101011),
      .k4(32'b10111101010111101101101101111110),
      .k5(32'b00111101011000110001010101011111),
      .k6(32'b10111100100001110111010100001001),
      .k7(32'b00111101110100100110010110110000),
      .k8(32'b10111101101000001001111000111101),
      .k9(32'b10111101110111001100111011111010)
  ) CON2D_13(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100101010001001110000111),
      .k2(32'b10111101010000100110010011001011),
      .k3(32'b00111101100001101011000111100111),
      .k4(32'b10111100100101011001110010011101),
      .k5(32'b10111101111000001111100111111011),
      .k6(32'b10111101011111101010110000110001),
      .k7(32'b10111101011001110111010101010011),
      .k8(32'b00111101001001000110001101000111),
      .k9(32'b10111101100111101100101111011011)
  ) CON2D_14(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100110010000100000010110010),
      .k2(32'b10111101100011110000010111000111),
      .k3(32'b10111101101001011101100100100000),
      .k4(32'b10111100100001001110001111010110),
      .k5(32'b00111100010110000111011101100110),
      .k6(32'b00111100011010111110010000001111),
      .k7(32'b00111100110101111011001001011001),
      .k8(32'b10111101111001111110001011011010),
      .k9(32'b10111101101000111100000010100000)
  ) CON2D_15(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101001001011000101111111),
      .k2(32'b10111101001010000010111101100100),
      .k3(32'b00111101101010100011011011000000),
      .k4(32'b00111100111000101111100001110011),
      .k5(32'b10111101100111101001000000010100),
      .k6(32'b00111101111110000000110010010101),
      .k7(32'b00111101101001010011000111001101),
      .k8(32'b10111101001000000101110001111100),
      .k9(32'b00111100011101001011000111010000)
  ) CON2D_16(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[0][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100010000011011111100110010)
)   op1(
    .i_pipeline_layer4(i_CORE_IP1[0]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*1-1:DATA_WIDTH*0])
);

/// CON2D_2///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101010001010110011001111),
      .k2(32'b10111101000000001101001010111011),
      .k3(32'b10111101010000010100010001001011),
      .k4(32'b10111101110010110000010111110011),
      .k5(32'b00111101000111101010000000001010),
      .k6(32'b00111101101010101000110100011110),
      .k7(32'b00111100101010101100110110101101),
      .k8(32'b10111101010000100100100110111001),
      .k9(32'b00111101000010101111111011001100)
  ) CON2D_17(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101100011000010001000111),
      .k2(32'b00111101100100010111001100111000),
      .k3(32'b00111100000101011111101001101101),
      .k4(32'b00111101110000001101101010111101),
      .k5(32'b00111100101000010010001001011111),
      .k6(32'b10111101111111000100100110001011),
      .k7(32'b10111101101100111110011110011111),
      .k8(32'b10111101111001100000010001001010),
      .k9(32'b00111011110011001011110000100001)
  ) CON2D_18(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010011111011011101111101),
      .k2(32'b10111101100001110011010100010000),
      .k3(32'b00111100100000110110001111000111),
      .k4(32'b10111101000011000011111010001111),
      .k5(32'b10111010101010010001101110010011),
      .k6(32'b10111101100001010011100011110010),
      .k7(32'b00111100011001111011101010111100),
      .k8(32'b10111101111100100100011100010001),
      .k9(32'b10111101110000110100100001010110)
  ) CON2D_19(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011101001001110100110110),
      .k2(32'b10111100111110100111010001011110),
      .k3(32'b10111101110111000110110111101010),
      .k4(32'b10111101101101111010110101011010),
      .k5(32'b10111101110110100001011101011110),
      .k6(32'b00111101110001010110001100100010),
      .k7(32'b00111101111111101000100101101100),
      .k8(32'b10111101001000111110100111101001),
      .k9(32'b10111100100011001101100000010010)
  ) CON2D_20(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111100000100010001101111),
      .k2(32'b10111100110100100111011011011100),
      .k3(32'b00111100110100111110110011001010),
      .k4(32'b10111101100010100001011101011110),
      .k5(32'b10111101000011111101100101011001),
      .k6(32'b00111101011000000000101011110001),
      .k7(32'b10111100110011100101010000110100),
      .k8(32'b10111101000110111000100010101101),
      .k9(32'b10111101110000101111000001100001)
  ) CON2D_21(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101011011011111001110011),
      .k2(32'b10111011011111110111010010111001),
      .k3(32'b00111100000011011001010011010110),
      .k4(32'b00111101110101001100010000101110),
      .k5(32'b00111100100010111111110110100111),
      .k6(32'b00111101101110111001100011101111),
      .k7(32'b00111101100010001010100011110001),
      .k8(32'b10111100110111011010010011000010),
      .k9(32'b10111101111001001011011101010111)
  ) CON2D_22(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001010110011010001100000),
      .k2(32'b00111101011000101110110101111101),
      .k3(32'b10111101100101000000000111001101),
      .k4(32'b10111101101000111001011001101001),
      .k5(32'b00111101101000110000000001010101),
      .k6(32'b10111101010001011010000000101100),
      .k7(32'b00111011001001100101100000110111),
      .k8(32'b10111101000111011110000011110010),
      .k9(32'b00111101101010010100010001111110)
  ) CON2D_23(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100010001000111000000100),
      .k2(32'b00111101110011111101010100001100),
      .k3(32'b00111101101011100110010101111001),
      .k4(32'b00111011111011011011111011011010),
      .k5(32'b00111101110111000101000101110111),
      .k6(32'b10111100011100010011010100101100),
      .k7(32'b10111101110011001110000000110010),
      .k8(32'b00111101001001101110000101000001),
      .k9(32'b10111101100000001101001000000111)
  ) CON2D_24(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111111011100100111011),
      .k2(32'b00111101100100000100110111011100),
      .k3(32'b10111010100000011000110010000001),
      .k4(32'b00111101000001000000011000000111),
      .k5(32'b10111101110000110110101010000100),
      .k6(32'b10111100110101110110001100110011),
      .k7(32'b00111100101111110000000010100111),
      .k8(32'b10111101011101111101100010010010),
      .k9(32'b10111101001001100000101001001010)
  ) CON2D_25(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111101010010010011000000),
      .k2(32'b00111100110000010010001010100100),
      .k3(32'b00111101100000010101111100110100),
      .k4(32'b10111101011101000010010110100001),
      .k5(32'b00111101111001011000100001100110),
      .k6(32'b10111101011010100011011110000110),
      .k7(32'b10111101001010000011101100111100),
      .k8(32'b00111101100010100110011111011010),
      .k9(32'b00111101111100110001111110010000)
  ) CON2D_26(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011000010111111111101),
      .k2(32'b10111100110000011111101101001010),
      .k3(32'b00111101010101010011111001001011),
      .k4(32'b10111101101001100011101101010100),
      .k5(32'b00111100110100110001111010010010),
      .k6(32'b10111101000000110010010010111001),
      .k7(32'b10111101100010110110010001111110),
      .k8(32'b00111100101111111110101011110100),
      .k9(32'b10111101101010100001100010100010)
  ) CON2D_27(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011101110010001111111101101),
      .k2(32'b10111101110101010010010000001110),
      .k3(32'b10111101001101000010110011010001),
      .k4(32'b10111100100101010011000111111001),
      .k5(32'b00111100101001101111100011000101),
      .k6(32'b10111110000000110001001001101011),
      .k7(32'b00111100111111110110010111100100),
      .k8(32'b00111010101000011100111111001000),
      .k9(32'b00111101000001000010110111111111)
  ) CON2D_28(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100001100000010110010001),
      .k2(32'b10111101001010111010100011010000),
      .k3(32'b10111011111101001100001100110110),
      .k4(32'b00111011111101110001010001100011),
      .k5(32'b00111100101000101110110011000000),
      .k6(32'b00111101111010110001110101001010),
      .k7(32'b10111100010101110110011011010011),
      .k8(32'b00111101100010011110110001101011),
      .k9(32'b00111101100110100111001011111000)
  ) CON2D_29(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111000010011011101010010),
      .k2(32'b00111100011100100101000011100111),
      .k3(32'b00111101001101000100011000111010),
      .k4(32'b10111101010101000101110010110011),
      .k5(32'b00111101100001011110111000010110),
      .k6(32'b10111011011100100100110001110011),
      .k7(32'b10111101011101101111010001001001),
      .k8(32'b10111101110010111000011000101100),
      .k9(32'b00111110000000101100000011010110)
  ) CON2D_30(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100100011101011100000111),
      .k2(32'b00111101110000010110010000000101),
      .k3(32'b10111100110011110101111111010100),
      .k4(32'b00111101001101101111111000001110),
      .k5(32'b00111101110010101100111000110110),
      .k6(32'b10111010010010010100001110110011),
      .k7(32'b10111101100001011010001010010101),
      .k8(32'b00111101111010001110111011100111),
      .k9(32'b00111101100000101010111001101011)
  ) CON2D_31(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100000111011010010100011),
      .k2(32'b10111100011011111010010111001000),
      .k3(32'b10111101100111000001111100011111),
      .k4(32'b00111101101100111100000111000111),
      .k5(32'b10111100101011011111111001100010),
      .k6(32'b10111100010111010100101000010010),
      .k7(32'b10111100001001000100100011001101),
      .k8(32'b10111010010110110010000011010011),
      .k9(32'b00111100001101010110100000001000)
  ) CON2D_32(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[1][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111001100001111100011010100101)
)   op2(
    .i_pipeline_layer4(i_CORE_IP1[1]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*2-1:DATA_WIDTH*1])
);

/// CON2D_3///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111111000101001010010000),
      .k2(32'b10111101100111001000011010000000),
      .k3(32'b00111101101000000111011100011100),
      .k4(32'b10111100001111111011101100111010),
      .k5(32'b10111100011010010110010000011101),
      .k6(32'b10111100110011111100110100100010),
      .k7(32'b10111101000110101100100001001001),
      .k8(32'b10111101110111000001011011011110),
      .k9(32'b00111101110001101110000101111101)
  ) CON2D_33(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011100110110100010110110001),
      .k2(32'b00111101011011011111111001100010),
      .k3(32'b00111101101010011100011100000000),
      .k4(32'b10111101001001000111101101000001),
      .k5(32'b10111101010010100001100100000101),
      .k6(32'b00111011100100101001100001001100),
      .k7(32'b10111101101011011111101100011010),
      .k8(32'b10111011110011010111001110110110),
      .k9(32'b10111101011000110011111111111101)
  ) CON2D_34(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000111101100111111011111),
      .k2(32'b10111101000101101001001111001001),
      .k3(32'b00111101100000010001010000100010),
      .k4(32'b00111100110011100100010110110110),
      .k5(32'b10111101110001110011000101111101),
      .k6(32'b10111101111000000100001011011110),
      .k7(32'b10111101000000101010011101001011),
      .k8(32'b10111101000010000000110110011010),
      .k9(32'b00111101001111000101110001011001)
  ) CON2D_35(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000111100001110100000000),
      .k2(32'b00111100110011100011000010110100),
      .k3(32'b00111101111100010101101100001011),
      .k4(32'b00111101011100011101010110010111),
      .k5(32'b00111011111010101101101000111101),
      .k6(32'b00111101111010111100101011011101),
      .k7(32'b00111100111000011101000101111101),
      .k8(32'b00111101110100001100001110001111),
      .k9(32'b10111101101101011000101001110000)
  ) CON2D_36(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111100111100000110011000),
      .k2(32'b10111100010000011000000101010110),
      .k3(32'b00111101100011111101100001111111),
      .k4(32'b10111101001000111101001110100111),
      .k5(32'b10111101101110000001010001110010),
      .k6(32'b00111101000000110011100111100111),
      .k7(32'b10111101101100101100101011000000),
      .k8(32'b10111101010010100110011000001101),
      .k9(32'b10111101001001110000101011010001)
  ) CON2D_37(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101111011000100010010100),
      .k2(32'b10111101000001100010001100010101),
      .k3(32'b00111101101100111111111110000000),
      .k4(32'b00111101100011010010101010100110),
      .k5(32'b00111101101001110010000101101110),
      .k6(32'b10111101010111111101110111001000),
      .k7(32'b10111101110101110111110101001110),
      .k8(32'b10111100110000001110010100000110),
      .k9(32'b10111011010010001010001111101001)
  ) CON2D_38(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111000010101001101000),
      .k2(32'b10111101110000100100110001101100),
      .k3(32'b10111100110100111011010101001000),
      .k4(32'b10111101000001001000111010000110),
      .k5(32'b10111101101101000010000101010010),
      .k6(32'b00111101000000011001010010011011),
      .k7(32'b00111110000010011001111011001001),
      .k8(32'b00111101101100100111110001100001),
      .k9(32'b00111101101001001011010101010011)
  ) CON2D_39(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011000001011011110010110),
      .k2(32'b10111101010011110111011001001111),
      .k3(32'b10111101100010001011000011011101),
      .k4(32'b00111101110001011100100010010010),
      .k5(32'b10111101101101111101100001111001),
      .k6(32'b00111101100000101111111100101000),
      .k7(32'b00111101101101000110000010010110),
      .k8(32'b00111101100101001111110011011000),
      .k9(32'b10111101000100110101000101010110)
  ) CON2D_40(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001101101101111001001011),
      .k2(32'b00111101101011100010111011011100),
      .k3(32'b00111101000010000101011111001000),
      .k4(32'b00111100000000000011111100111101),
      .k5(32'b10111101110001000010001101110000),
      .k6(32'b00111101001111100100111100010000),
      .k7(32'b00111101110101110100111010100010),
      .k8(32'b10111100111011100000000001100110),
      .k9(32'b00111101011011011101101100101110)
  ) CON2D_41(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111001000100011010111011),
      .k2(32'b10111101101000100001100101001111),
      .k3(32'b10111011001100111100101101001100),
      .k4(32'b00111101010110100001001101001000),
      .k5(32'b10111101101000100111000101111110),
      .k6(32'b10111101000000100011101010100110),
      .k7(32'b10111101011000100100010111010011),
      .k8(32'b10111101101011101110101101001101),
      .k9(32'b00111101000001111001100101011110)
  ) CON2D_42(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001100111110000001111),
      .k2(32'b10111101101100001001001011010101),
      .k3(32'b10111100110111101010000011111100),
      .k4(32'b00111101110001101010111111010010),
      .k5(32'b10111101101110100011011110101111),
      .k6(32'b10111100111010011010001011110010),
      .k7(32'b00111101101000001110010100011011),
      .k8(32'b10111101100100011101001001111001),
      .k9(32'b10111101111011001010011111111010)
  ) CON2D_43(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110100001010001010110011),
      .k2(32'b10111101100111100111111100101111),
      .k3(32'b00111101101110111100101111001110),
      .k4(32'b10111101000000001110000101011010),
      .k5(32'b00111101111111011111111010110000),
      .k6(32'b00111101001000001000010111000111),
      .k7(32'b00111101111110100001010111110001),
      .k8(32'b00111101001001100000011111100110),
      .k9(32'b00111101111011101011000000100101)
  ) CON2D_44(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011011001110010001010110),
      .k2(32'b10111100110001000010100001110000),
      .k3(32'b00111101111010011010010011111100),
      .k4(32'b00111101101011101110110110111001),
      .k5(32'b00111101110111001011001111100110),
      .k6(32'b10111101010011011101100110001001),
      .k7(32'b10111101100011111010111100110111),
      .k8(32'b00111101110111001101110010001110),
      .k9(32'b00111100001000111111110110011110)
  ) CON2D_45(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110001001010000101101011),
      .k2(32'b00111100011001001110111011000010),
      .k3(32'b00111100100101100010111000000010),
      .k4(32'b00111101110000111110101110010011),
      .k5(32'b10111011101100110010110110100010),
      .k6(32'b10111101101011001010111101011100),
      .k7(32'b10111100101101000010001000110000),
      .k8(32'b00111101100111001000000010101010),
      .k9(32'b10111101001001111010101110011110)
  ) CON2D_46(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011110110110110110110),
      .k2(32'b10111101101100001010001111110001),
      .k3(32'b10111110000000101011010111101100),
      .k4(32'b00111011001100011101100001010001),
      .k5(32'b10111100110000001100000001010011),
      .k6(32'b00111101001001000011001101001111),
      .k7(32'b00111011111101011100110000111001),
      .k8(32'b10111101101011111010010000100111),
      .k9(32'b10111101111001100000100001010011)
  ) CON2D_47(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101111100000000000011100),
      .k2(32'b00111101110000101100001101001000),
      .k3(32'b10111101110001111111001010101111),
      .k4(32'b10111100100100011000000100011011),
      .k5(32'b10111100100001101000000001111100),
      .k6(32'b00111100011010110101001111000010),
      .k7(32'b10111101011001100001100111101100),
      .k8(32'b00111011101110100011000000001000),
      .k9(32'b10111101010101100101100010101101)
  ) CON2D_48(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[2][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100100010110111001100100101)
)   op3(
    .i_pipeline_layer4(i_CORE_IP1[2]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*3-1:DATA_WIDTH*2])
);

/// CON2D_4///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100110101000100111011001110),
      .k2(32'b00111100101000000100101101110010),
      .k3(32'b10111101010001000111101111001110),
      .k4(32'b10111101011011000011101010111010),
      .k5(32'b10111101000000100110011001001110),
      .k6(32'b00111101001001111111011000011110),
      .k7(32'b00111101100010011111000000001001),
      .k8(32'b10111101011001000001010010001100),
      .k9(32'b00111101111000011000110010000100)
  ) CON2D_49(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000001111010001001000111),
      .k2(32'b10111100111001001000000100010101),
      .k3(32'b00111100101011000100010111101111),
      .k4(32'b00111101110111011100010010000000),
      .k5(32'b00111110000011011100011010010110),
      .k6(32'b10111100110110101110000001011111),
      .k7(32'b00111100000111000011101000111110),
      .k8(32'b00111101010100000011010011001110),
      .k9(32'b10111010101111101011011110110110)
  ) CON2D_50(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010011011011001101000111),
      .k2(32'b00111100111100011110100001010001),
      .k3(32'b00111101110111011100110110000001),
      .k4(32'b10111100110111101110000111110111),
      .k5(32'b00111100010110011001110110110101),
      .k6(32'b10111101100101001000011100011101),
      .k7(32'b00111100111110001000011101100110),
      .k8(32'b10111100001101100010110111000001),
      .k9(32'b00111101011010010111001100011010)
  ) CON2D_51(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101000010110000101100010),
      .k2(32'b10111101110110010000101110111110),
      .k3(32'b10111100101100010000111101011111),
      .k4(32'b00111100011010010110110111000000),
      .k5(32'b10111101001101001111101111111011),
      .k6(32'b10111100110101100111001110110110),
      .k7(32'b00111101100100110001011111111000),
      .k8(32'b00111101101110011111010001101011),
      .k9(32'b00111101101101001010101010100111)
  ) CON2D_52(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101000001100110010000001),
      .k2(32'b10111101001101010011101111001101),
      .k3(32'b00111101101101001000101011000001),
      .k4(32'b10111101010111000000101000010011),
      .k5(32'b10111011111110011010110111001001),
      .k6(32'b00111101110010100101010100010000),
      .k7(32'b00111100010010111001010110001111),
      .k8(32'b00111101000111111010001111010001),
      .k9(32'b00111101111011100010001101100001)
  ) CON2D_53(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010010011111111010100011),
      .k2(32'b10111100101001100001100101110000),
      .k3(32'b10111100101110100010000011111110),
      .k4(32'b10111101110111001010011010000000),
      .k5(32'b10111100011011000110110111100001),
      .k6(32'b10111101110000101010101010110100),
      .k7(32'b10111100000101100010010000000111),
      .k8(32'b00111101110011001011101110100001),
      .k9(32'b10111101000011111000011000010101)
  ) CON2D_54(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000001011001101010001010),
      .k2(32'b10111101011011001110001110000010),
      .k3(32'b10111101001111110001010110010001),
      .k4(32'b00111101111000101100100100101010),
      .k5(32'b00111100000110000101001100110001),
      .k6(32'b00111011111101100011100011101111),
      .k7(32'b00111101100100000001011011001010),
      .k8(32'b00111101000010101101000011110011),
      .k9(32'b00111101110001111101100101101110)
  ) CON2D_55(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101001101101010100110111),
      .k2(32'b10111101010010000010010010001100),
      .k3(32'b00111100110101001111001001110000),
      .k4(32'b10111101101010010000110000101100),
      .k5(32'b00111100011001100100100010011001),
      .k6(32'b00111101110011111101100000110010),
      .k7(32'b00111101100110110111110110110000),
      .k8(32'b10111101000000111010000110111000),
      .k9(32'b10111101101000011110101100111101)
  ) CON2D_56(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111010111100010011011110),
      .k2(32'b10111101000000001001010010111101),
      .k3(32'b10111001100110011001001000000010),
      .k4(32'b10111101110000110010000001000101),
      .k5(32'b10111101001001011011001101111110),
      .k6(32'b00111100010001111100001001101101),
      .k7(32'b10111101011101011110100010100111),
      .k8(32'b00111100100011110100101010100000),
      .k9(32'b00111101111011010011111101111000)
  ) CON2D_57(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100111010111000011100101),
      .k2(32'b00111101110101001011010011101111),
      .k3(32'b00111100110010001101101001100100),
      .k4(32'b00111101100100100001101010111111),
      .k5(32'b00111100100010001011110101001001),
      .k6(32'b10111100011011000000011100100101),
      .k7(32'b10111100100110001011000001001000),
      .k8(32'b00111101001101001111000101000000),
      .k9(32'b10111101010101000111011100001110)
  ) CON2D_58(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110111001111010100101101),
      .k2(32'b00111101100000011100110111001101),
      .k3(32'b10111101011011110001110110101110),
      .k4(32'b00111011111011110101011111001011),
      .k5(32'b10111101000101111011011101100111),
      .k6(32'b10111101100000110010100000000011),
      .k7(32'b10111101101100001110011111111100),
      .k8(32'b10111100101111001111000100110001),
      .k9(32'b10111011100011000110110000101100)
  ) CON2D_59(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011100001011110000000100),
      .k2(32'b10111101100000011010011010011111),
      .k3(32'b00111101011010101110110011010111),
      .k4(32'b10111010101001010101010000011111),
      .k5(32'b00111100110111111001100111011000),
      .k6(32'b00111101100100111000111010010000),
      .k7(32'b00111101100111100010000000110000),
      .k8(32'b00111100010100111101100001011010),
      .k9(32'b10111101011100001100111010101100)
  ) CON2D_60(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100001010011111111111111),
      .k2(32'b10111011111101100101011110010110),
      .k3(32'b10111101101100000010110110001000),
      .k4(32'b00111101010110001011101111111100),
      .k5(32'b10111100110010000001110111011000),
      .k6(32'b00111101100011110100111000100011),
      .k7(32'b10111101100110010111000000111111),
      .k8(32'b10111101111011000001111101000101),
      .k9(32'b10111101100001110100100110110110)
  ) CON2D_61(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110100101111101011001),
      .k2(32'b00111101111000100101101110110001),
      .k3(32'b00111101101001110101000011010010),
      .k4(32'b10111101101101011101110100001010),
      .k5(32'b10111101111011100100010001100011),
      .k6(32'b00111101100011011111111010000000),
      .k7(32'b00111100110100101101000011001101),
      .k8(32'b00111100001011110001010110001011),
      .k9(32'b00111101110010011111110101011010)
  ) CON2D_62(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110000001011001100101),
      .k2(32'b10111011011010101010001010001010),
      .k3(32'b10111101000001110100011001110001),
      .k4(32'b10111101000001101001110000000100),
      .k5(32'b00111100010010111110100011100010),
      .k6(32'b10111101111000000010010111111111),
      .k7(32'b10111101010011101111010101110101),
      .k8(32'b00111101011101101110100001000011),
      .k9(32'b00111101001000110101010001000111)
  ) CON2D_63(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001000010111011110001010),
      .k2(32'b00111101001110010100000111001101),
      .k3(32'b10111010001101011110001100100011),
      .k4(32'b00111101110010110100111000010111),
      .k5(32'b10111011000010010111101010111011),
      .k6(32'b10111100100011111010000100000100),
      .k7(32'b10111010001110011110000011011010),
      .k8(32'b00111100000001001011011011100101),
      .k9(32'b00111101111100000100000001100001)
  ) CON2D_64(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[3][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100101000100110010111100111)
)   op4(
    .i_pipeline_layer4(i_CORE_IP1[3]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*4-1:DATA_WIDTH*3])
);

/// CON2D_5///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011001010001011100010000),
      .k2(32'b00111000111110000110011000001101),
      .k3(32'b00111101101010111000000001101100),
      .k4(32'b00111100111001001001000011101000),
      .k5(32'b10111101011011100101111111101111),
      .k6(32'b00111100000100110011111101101110),
      .k7(32'b10111101100110001111111100111010),
      .k8(32'b00111101100101111011001101000110),
      .k9(32'b10111011001110010000100000100110)
  ) CON2D_65(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001011111001101011110011),
      .k2(32'b10111101110101110001111110000011),
      .k3(32'b00111101101011101011100110111010),
      .k4(32'b10111100110101101100001000001100),
      .k5(32'b10111101110001010000011110110100),
      .k6(32'b10111100001111101000111010110011),
      .k7(32'b00111101001101100100101111001000),
      .k8(32'b10111100110101110000001010100001),
      .k9(32'b10111101111000001011001011110110)
  ) CON2D_66(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101001001011100011011001),
      .k2(32'b00111100111010000011101010100110),
      .k3(32'b10111101100011111000110011001011),
      .k4(32'b00111101000111001111111001110110),
      .k5(32'b00111101101111001110111010100110),
      .k6(32'b00111101001000101110011111010001),
      .k7(32'b10111101111011110101100101010100),
      .k8(32'b00111100110000011100100111011001),
      .k9(32'b10111101100100111001000010110110)
  ) CON2D_67(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111001000010010100001000),
      .k2(32'b10111101110000000000110010001001),
      .k3(32'b00111101101010011000110110001010),
      .k4(32'b10111101000011101110001101110111),
      .k5(32'b00111101001000001000101000000001),
      .k6(32'b00111101111010111001100001010010),
      .k7(32'b00111101001101101100110011100011),
      .k8(32'b10111101101010010110011110100010),
      .k9(32'b00111101001010110101100111000101)
  ) CON2D_68(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110010110111100110010),
      .k2(32'b00111101100111010111110001010100),
      .k3(32'b00111101101110000001110001010011),
      .k4(32'b00111100100010111110100001100111),
      .k5(32'b00111101001110001011111100100100),
      .k6(32'b00111011101111101010000010010010),
      .k7(32'b10111100011010110100101001110011),
      .k8(32'b10111101111110000001011101000110),
      .k9(32'b10111101101011100011101100001001)
  ) CON2D_69(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010111010010010001011),
      .k2(32'b10111100101001001011100000101111),
      .k3(32'b10111101101000110101110001001110),
      .k4(32'b10111101011110010001100111010100),
      .k5(32'b00111101111010001100110111110001),
      .k6(32'b00111100110001010110001111111010),
      .k7(32'b00111100111010100010000100111100),
      .k8(32'b00111101110001100100001110100011),
      .k9(32'b00111100101101101000110111111010)
  ) CON2D_70(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110101000111011000000111),
      .k2(32'b00111101110101110110101101101010),
      .k3(32'b00111101001001101001111101001000),
      .k4(32'b00111100111101110101110110000000),
      .k5(32'b00111100100110000011001100011100),
      .k6(32'b10111101010110011101110001111100),
      .k7(32'b10111101100010101100111111110110),
      .k8(32'b00111101111000010101001010010111),
      .k9(32'b10111101001000010010101100111001)
  ) CON2D_71(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011010000100010110010000),
      .k2(32'b00111101010110001001001010101010),
      .k3(32'b00111101101101101010001010000001),
      .k4(32'b10111101000111000100100100110010),
      .k5(32'b00111101000001100101101111110001),
      .k6(32'b00111101110100111111111100001001),
      .k7(32'b00111101010000111000010100011111),
      .k8(32'b00111101111100100001111011111101),
      .k9(32'b10111101110111110100100011101010)
  ) CON2D_72(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010000011100000101001100),
      .k2(32'b00111100010010011100110111001101),
      .k3(32'b00111101000111101010100000010000),
      .k4(32'b10111101000000100100010100000000),
      .k5(32'b00111101011001010111111010111011),
      .k6(32'b00111100000001100110011101101011),
      .k7(32'b00111101101100101000010100100000),
      .k8(32'b10111101111111000011000111111101),
      .k9(32'b00111100110111111001000101000001)
  ) CON2D_73(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100100000001100100011010),
      .k2(32'b10111100011101101000011111000011),
      .k3(32'b10111101000100001010001100010110),
      .k4(32'b10111101101000001110110010011010),
      .k5(32'b10111101000000111010110011111101),
      .k6(32'b00111101010000100000001001111111),
      .k7(32'b00111101000010000000011000111001),
      .k8(32'b00111100111100011111010011101100),
      .k9(32'b00111101011011001101100010000101)
  ) CON2D_74(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100100001101011100010),
      .k2(32'b00111101110001111010001101011100),
      .k3(32'b00111101011100101101001110110111),
      .k4(32'b00111101111001000000101101000010),
      .k5(32'b00111011100101010011010010010100),
      .k6(32'b10111101011011001011100101100011),
      .k7(32'b00111101101111000100011010000111),
      .k8(32'b10111101001101000000111111001111),
      .k9(32'b10111101101011000011100101100110)
  ) CON2D_75(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110011001011111111000101),
      .k2(32'b10111011100001011100101011111110),
      .k3(32'b10111100110010011010000110100001),
      .k4(32'b10111011100011111000101000100100),
      .k5(32'b00111100010011110001000000100100),
      .k6(32'b00111101110010010111111001110101),
      .k7(32'b10111100111101110001111011110011),
      .k8(32'b10111101000011010110110111001110),
      .k9(32'b00111101001011000110111110001111)
  ) CON2D_76(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100011011110001011110),
      .k2(32'b00111101001111110101101111111011),
      .k3(32'b10111101000100101101111000001110),
      .k4(32'b10111100110000111010010111000001),
      .k5(32'b10111101001100101111111100110110),
      .k6(32'b10111101111001110101001000001000),
      .k7(32'b00111101110001001001000010110011),
      .k8(32'b10111100100001011100101001110011),
      .k9(32'b00111101011011101111101110110101)
  ) CON2D_77(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100100011000110010101111),
      .k2(32'b10111101010111000011000110110111),
      .k3(32'b10111101100001100001010010001110),
      .k4(32'b10111101001110011010001110010111),
      .k5(32'b00111101110011001100010010011000),
      .k6(32'b00111101000111101000001011101011),
      .k7(32'b00111100010011111011010110000011),
      .k8(32'b10111101000010100000111100011010),
      .k9(32'b10111100111011110111101111001000)
  ) CON2D_78(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100010101101010000010111),
      .k2(32'b00111100111100011101111111011010),
      .k3(32'b10111101111110101011111001011110),
      .k4(32'b00111101111101111000111000000000),
      .k5(32'b10111011111101001111100110001110),
      .k6(32'b10111101101111000101110100111011),
      .k7(32'b10111101100111001110111001100100),
      .k8(32'b00111101100001100010001011101001),
      .k9(32'b10111101000011001011010100100011)
  ) CON2D_79(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010011111011110001110110),
      .k2(32'b00111101000010001111111110111010),
      .k3(32'b00111101110101100010100011100111),
      .k4(32'b10111101101010111001001101111011),
      .k5(32'b10111101111100100100001010111101),
      .k6(32'b00111011100010000001011000111100),
      .k7(32'b10111101100101011101111110110000),
      .k8(32'b10111101101101011001111101101111),
      .k9(32'b10111100001100111001100000101110)
  ) CON2D_80(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[4][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111100000010000011100101010011)
)   op5(
    .i_pipeline_layer4(i_CORE_IP1[4]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*5-1:DATA_WIDTH*4])
);

/// CON2D_6///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101110001011010010101010),
      .k2(32'b00111101101011000110101110000101),
      .k3(32'b00111101111011011010110101100000),
      .k4(32'b10111101001100001010100110011011),
      .k5(32'b10111100001011111111011111101010),
      .k6(32'b00111101110110101101000000100011),
      .k7(32'b10111101100111010011111011101110),
      .k8(32'b10111101110000011000000000100010),
      .k9(32'b00111101110000000110111000110001)
  ) CON2D_81(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111001000100111110001110),
      .k2(32'b10111101101011111111100101001110),
      .k3(32'b10111101101111101100100000000001),
      .k4(32'b00111101110011111110101000000100),
      .k5(32'b00111100100010100011101001010001),
      .k6(32'b00111101010111111101001101000010),
      .k7(32'b00111100101011110100110101010101),
      .k8(32'b10111001111110101001011101011100),
      .k9(32'b10111101110011011001010011111010)
  ) CON2D_82(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111100101000111001010010),
      .k2(32'b00111100001001111001101000011101),
      .k3(32'b10111100000111000101000011100101),
      .k4(32'b10111101100101001001110010011011),
      .k5(32'b10111101100100110100111111011000),
      .k6(32'b10111100101000011111011000000000),
      .k7(32'b10111101011000100010000000100101),
      .k8(32'b10111101100100000000101100101011),
      .k9(32'b10111101010001101110000101000101)
  ) CON2D_83(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010111000011000010111),
      .k2(32'b00111101101101100011010101000111),
      .k3(32'b10111101111001011111111011100011),
      .k4(32'b10111101110000101011001101100001),
      .k5(32'b10111100100000000101100010011011),
      .k6(32'b00111100111011000101100001001111),
      .k7(32'b10111101000001111101100111110001),
      .k8(32'b10111101100001111100110101111011),
      .k9(32'b00111101000011011100111101010011)
  ) CON2D_84(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001001101111111001111100),
      .k2(32'b00111101100011010110101001101010),
      .k3(32'b10111101110100101100010000111010),
      .k4(32'b10111101010001100011110000010111),
      .k5(32'b10111101001000111001101011110010),
      .k6(32'b00111101100111110111100011000010),
      .k7(32'b00111101101101001011001011011111),
      .k8(32'b10111101111101000001100110000000),
      .k9(32'b00111101010101001010010101001101)
  ) CON2D_85(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100000011000110011001000),
      .k2(32'b10111011101110101010000000001110),
      .k3(32'b10111100111110111001000111101011),
      .k4(32'b00111100110101110001011011101100),
      .k5(32'b10111101100010001010011110000101),
      .k6(32'b10111101000011101101000110111110),
      .k7(32'b10111101001011101000110000001010),
      .k8(32'b10111101111110101110111100101010),
      .k9(32'b10111100111010010101001001001111)
  ) CON2D_86(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110000010000010011110110),
      .k2(32'b10111101100100001100010001110000),
      .k3(32'b00111011111001011110101010101100),
      .k4(32'b10111100010110011011010011101101),
      .k5(32'b10111101111010000010010111000101),
      .k6(32'b10111101001100111000100100101101),
      .k7(32'b00111101001101010110100110100110),
      .k8(32'b00111101001100111001000111011101),
      .k9(32'b00111100001100110001010010100101)
  ) CON2D_87(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011110011111011110111000110),
      .k2(32'b00111100000101100101010101001000),
      .k3(32'b00111101100001000010001110000110),
      .k4(32'b00111101100110101000101100001101),
      .k5(32'b00111101110100110111000000000110),
      .k6(32'b10111100010010011011001111100100),
      .k7(32'b00111100000000110000100100011101),
      .k8(32'b10111100100101000111001100101011),
      .k9(32'b00111100110101001011001010010110)
  ) CON2D_88(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100010111110000110001000),
      .k2(32'b10111100100011110111011001100011),
      .k3(32'b00111100100101011001010000110001),
      .k4(32'b10111101111111100001001111110011),
      .k5(32'b00111100110111111011000011010101),
      .k6(32'b10111101110100001001011100010000),
      .k7(32'b00111010110000000010010111010110),
      .k8(32'b10111101101011101011001111000010),
      .k9(32'b10111101110101100001101111110111)
  ) CON2D_89(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111000000011100100010),
      .k2(32'b10111101100110101010100100110111),
      .k3(32'b00111101101101101000001110010110),
      .k4(32'b00111101000101101101011111110010),
      .k5(32'b10111101010001000110010101010011),
      .k6(32'b10111100101110101111011100111101),
      .k7(32'b10111101000011100110101000110101),
      .k8(32'b10111101000111010100000101011110),
      .k9(32'b00111101011011100110000010011100)
  ) CON2D_90(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100101100101100101010001),
      .k2(32'b00111101101000000000110111011111),
      .k3(32'b10111101110001010000011110000100),
      .k4(32'b10111011001100101001110110001011),
      .k5(32'b00111101110111000110101101111001),
      .k6(32'b10111101000100111001110000001000),
      .k7(32'b10111101001101100011100101001111),
      .k8(32'b00111101101110111001111010001010),
      .k9(32'b00111101110110011010000011001111)
  ) CON2D_91(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011101010101011000010101),
      .k2(32'b10111100111000011000011100011011),
      .k3(32'b00111101010001101011001011011111),
      .k4(32'b10111011110000101100011101001001),
      .k5(32'b10111101101010100000001011001011),
      .k6(32'b10111110000100010000100100101001),
      .k7(32'b00111101101010000110010001011110),
      .k8(32'b10111101110101011011011110000111),
      .k9(32'b10111110000111111100101111011010)
  ) CON2D_92(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011101010011100100010000101),
      .k2(32'b10111101010001001001101010101010),
      .k3(32'b10111101100001101101101010111000),
      .k4(32'b10111100100010001000011101110111),
      .k5(32'b00111101110110110110110000101011),
      .k6(32'b10111100110111111000101011111101),
      .k7(32'b10111101110101100010001011010110),
      .k8(32'b10111100110000010111110010001110),
      .k9(32'b10111101100011001010101110100111)
  ) CON2D_93(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111001010111100001110101),
      .k2(32'b00111100101011011101000000010011),
      .k3(32'b00111101011010100111011001000000),
      .k4(32'b00111101010100000100110111100011),
      .k5(32'b00111100111001100101101111100111),
      .k6(32'b10111101000000110101111010000000),
      .k7(32'b00111101101110011001011001100111),
      .k8(32'b00111101001110111000100011100011),
      .k9(32'b10111101010110000000010010001111)
  ) CON2D_94(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100000010000111111000011101),
      .k2(32'b10111101100111001100010000011100),
      .k3(32'b00111011101111011100100110000000),
      .k4(32'b10111101101011010111001011001101),
      .k5(32'b00111110000011000110110110000010),
      .k6(32'b00111100111010110001011000000001),
      .k7(32'b00111101001101011011101100111100),
      .k8(32'b00111110000100000110010110011100),
      .k9(32'b10111101100100010010010010101001)
  ) CON2D_95(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100101000111110000011),
      .k2(32'b00111101110110101001011011011011),
      .k3(32'b00111101011111001010011100110010),
      .k4(32'b00111101101010001100111001101001),
      .k5(32'b00111101110001011011101101101011),
      .k6(32'b10111101111000101101010101010110),
      .k7(32'b10111101011000101011110001000000),
      .k8(32'b00111101010000000001010101010010),
      .k9(32'b10111100010100111011110000010001)
  ) CON2D_96(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[5][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011100111100011100011001101)
)   op6(
    .i_pipeline_layer4(i_CORE_IP1[5]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*6-1:DATA_WIDTH*5])
);

/// CON2D_7///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110101110111100001010),
      .k2(32'b10111101101000011001111011110110),
      .k3(32'b00111101000111001101110000101100),
      .k4(32'b00111101001011001111100000110001),
      .k5(32'b00111101010011011000100110110001),
      .k6(32'b10111010001111001000111000101111),
      .k7(32'b00111100100100011011000010011011),
      .k8(32'b00111101110111110110111111100011),
      .k9(32'b10111101100011110001110111110001)
  ) CON2D_97(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100101100001000011111100),
      .k2(32'b10111101101010001011010110010000),
      .k3(32'b00111100001001000100011000111100),
      .k4(32'b10111100100011011011010100100011),
      .k5(32'b00111101011011010101001011110001),
      .k6(32'b10111011110000100010011011110101),
      .k7(32'b10111101101011000111100100010111),
      .k8(32'b10111100110101011011101000000110),
      .k9(32'b10111101101101100011001001010110)
  ) CON2D_98(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010100110100101011001000),
      .k2(32'b00111101001110011110100001100001),
      .k3(32'b10111101100011001100100110010001),
      .k4(32'b00111101101010001111011101011000),
      .k5(32'b00111101101111010001001011010011),
      .k6(32'b00111101010110110000011101100111),
      .k7(32'b10111011110110110111001101010101),
      .k8(32'b10111101100010010000110001010110),
      .k9(32'b00111101011111111100101011011001)
  ) CON2D_99(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100010011110100110000000),
      .k2(32'b10111101010011001110111011110100),
      .k3(32'b10111011101010100110010110101000),
      .k4(32'b00111100010110000111111011000100),
      .k5(32'b00111101101011010110111111001000),
      .k6(32'b00111101110101000101101111110011),
      .k7(32'b10111101001101000000000111100001),
      .k8(32'b00111101101010111110101100001001),
      .k9(32'b00111100110111100100001001011110)
  ) CON2D_100(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011101011000101100111001),
      .k2(32'b00111101100011000110111101100000),
      .k3(32'b00111101110001110111101001001111),
      .k4(32'b00111100001101010111001110010011),
      .k5(32'b00111100110110111010110110100111),
      .k6(32'b00111101110000111111011101100111),
      .k7(32'b00111101111001101100110101101011),
      .k8(32'b10111101110010100111110111110111),
      .k9(32'b10111101110001110101100110000111)
  ) CON2D_101(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011101011110111011110010),
      .k2(32'b00111101100111011000110010100010),
      .k3(32'b10111100011111110001111110101010),
      .k4(32'b00111101111000111111110110100000),
      .k5(32'b10111101100111111000000000101000),
      .k6(32'b00111101010111001110100000110100),
      .k7(32'b00111101101101100011110010101000),
      .k8(32'b00111100111000010100100011000011),
      .k9(32'b00111101101010110011101110001010)
  ) CON2D_102(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001110001111111001000111),
      .k2(32'b00111101101110000010000110100010),
      .k3(32'b00111101110000100011000101111111),
      .k4(32'b00111100010001110010010001001111),
      .k5(32'b10111100110001101101011110111001),
      .k6(32'b10111101100110101000100001011011),
      .k7(32'b10111101001001000101000001110111),
      .k8(32'b10111100111101011110110011100001),
      .k9(32'b00111101001011010101110101110110)
  ) CON2D_103(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101000011110101011101000),
      .k2(32'b00111101001001100011010111011000),
      .k3(32'b10111101100111001100110100010101),
      .k4(32'b10111101011001011011100101001011),
      .k5(32'b00111101000011101000101111110010),
      .k6(32'b00111011111100000011111001011001),
      .k7(32'b00111101111010001010000101100001),
      .k8(32'b10111101010000100101000111011111),
      .k9(32'b10111101000111101011101111100000)
  ) CON2D_104(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010111010011010110000111),
      .k2(32'b00111101100110011011011100100011),
      .k3(32'b10111101110001011100001011011100),
      .k4(32'b00111101100101001011100101010001),
      .k5(32'b10111101111001011111111011011010),
      .k6(32'b00111101110100011111000110111111),
      .k7(32'b00111101011011000011110011101001),
      .k8(32'b10111101111110010110000101001111),
      .k9(32'b00111100100101101001100101011110)
  ) CON2D_105(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110111001111110110000101),
      .k2(32'b10111101111011100101100101001111),
      .k3(32'b10111101101100100001110111100111),
      .k4(32'b00111101100100010110111101110001),
      .k5(32'b10111101110100100110001010011010),
      .k6(32'b10111100111010000000110111110101),
      .k7(32'b10111101010011001001000011100010),
      .k8(32'b10111101101100110110100000111001),
      .k9(32'b00111101011100100100101111001000)
  ) CON2D_106(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011110100011000111001000),
      .k2(32'b10111101100001110001010001011010),
      .k3(32'b10111101000011100000100101110111),
      .k4(32'b00111101100010010001010011001110),
      .k5(32'b00111101101100110011110010010111),
      .k6(32'b00111101100010011101110101000110),
      .k7(32'b10111100001000111111010100011010),
      .k8(32'b00111101001000000001001011110110),
      .k9(32'b00111101010110011100001110111100)
  ) CON2D_107(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111010111010010111001111111100),
      .k2(32'b00111101101000011111011011000110),
      .k3(32'b00111011001110100010111000111100),
      .k4(32'b00111101111001101110110101000110),
      .k5(32'b00111101011010111010110100100001),
      .k6(32'b10111100110101000000011010000100),
      .k7(32'b10111101111010110000111110110010),
      .k8(32'b00111101101100101111010111110111),
      .k9(32'b00111101110110101111101101000100)
  ) CON2D_108(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101111000110010111101100),
      .k2(32'b00111101011100101011100100001011),
      .k3(32'b10111101110110110101001111011001),
      .k4(32'b00111101100010000110110100100001),
      .k5(32'b10111010110010000111000100101011),
      .k6(32'b00111100000000001110100110100111),
      .k7(32'b00111101100101010000001101100000),
      .k8(32'b10111101010010000010010010000010),
      .k9(32'b10111101110111100011110001001000)
  ) CON2D_109(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001010101100011000111100),
      .k2(32'b10111101011001001010100001100000),
      .k3(32'b10111100100000101101101101101010),
      .k4(32'b10111101110011000100101110010101),
      .k5(32'b10111100010011010000001110101011),
      .k6(32'b00111101000011110010001110100101),
      .k7(32'b00111101100110110010111110101111),
      .k8(32'b00111101000111100110001101110011),
      .k9(32'b00111101100111100100010101010010)
  ) CON2D_110(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101010000011101001111010),
      .k2(32'b00111101101100010101011000001101),
      .k3(32'b10111101001010101011011000101110),
      .k4(32'b00111100011000000011101100110010),
      .k5(32'b00111100110110011000011001111110),
      .k6(32'b10111101101010010001110000000011),
      .k7(32'b00111101000000011111000011011001),
      .k8(32'b00111100001000001101011011000100),
      .k9(32'b00111101000011001101011001111100)
  ) CON2D_111(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111100001100010101010100),
      .k2(32'b00111101111110110111100011000010),
      .k3(32'b10111011110000010000010010111101),
      .k4(32'b10111100101010111111101001111100),
      .k5(32'b00111101100111101011000111011111),
      .k6(32'b10111101110101110111001010001001),
      .k7(32'b00111101100000000011011000001101),
      .k8(32'b10111101101000000101110010100100),
      .k9(32'b10111101010100101001101110010010)
  ) CON2D_112(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[6][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111010100100100110000000010010)
)   op7(
    .i_pipeline_layer4(i_CORE_IP1[6]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*7-1:DATA_WIDTH*6])
);

/// CON2D_8///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100101111011011001010001),
      .k2(32'b00111101110110111011010011101100),
      .k3(32'b00111101100010100001100010101000),
      .k4(32'b00111101111001111000111001001110),
      .k5(32'b10111101111010011100001001111101),
      .k6(32'b00111100110000011110110011110001),
      .k7(32'b10111100000011110100111000110011),
      .k8(32'b00111101100111101111100100101101),
      .k9(32'b00111100101011111010110011101110)
  ) CON2D_113(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011110001001001111101100),
      .k2(32'b00111101111000110000101000110101),
      .k3(32'b10111100101111000101101100001011),
      .k4(32'b10111101110010010110010101000100),
      .k5(32'b00111101010000001000111101011011),
      .k6(32'b00111101110101101110010011001111),
      .k7(32'b00111101001100110000001101010011),
      .k8(32'b10111101100011110001000111110001),
      .k9(32'b10111100101111110001100111100000)
  ) CON2D_114(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011000011100000011110101),
      .k2(32'b00111101100010101000010010111101),
      .k3(32'b00111011100111011011000000101110),
      .k4(32'b10111010000101111110011101010100),
      .k5(32'b00111101110001011111111011011000),
      .k6(32'b10111100101101010101111001100101),
      .k7(32'b00111101101101111011100000010111),
      .k8(32'b10111101101000001101100000111001),
      .k9(32'b10111101110101100111000000001101)
  ) CON2D_115(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010001101011001010000),
      .k2(32'b10111101101001100001110110011101),
      .k3(32'b00111101101001111010111001110101),
      .k4(32'b00111100001010110010101011111111),
      .k5(32'b10111101100100111110001100100101),
      .k6(32'b00111011100101101001011000000011),
      .k7(32'b00111101010101101101001101000111),
      .k8(32'b00111100011011110010000000011100),
      .k9(32'b00111100100101101000000001001000)
  ) CON2D_116(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010100001111010100011101),
      .k2(32'b00111101100111001100111101101001),
      .k3(32'b00111101001101100011101000101001),
      .k4(32'b10111101100111010111110011000110),
      .k5(32'b00111101110011000101011000001111),
      .k6(32'b00111101011001001000100001111011),
      .k7(32'b00111101110010010100000011000010),
      .k8(32'b10111101100100001011110100101010),
      .k9(32'b00111101100000110110000001111101)
  ) CON2D_117(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011010111010001000010),
      .k2(32'b00111100110010000000011111110101),
      .k3(32'b10111101110010101100001001010011),
      .k4(32'b10111100100100111011011011001011),
      .k5(32'b10111101110011100001000111000101),
      .k6(32'b00111101100110101011110101010110),
      .k7(32'b00111101010110110001011001100101),
      .k8(32'b10111101110111100011010011001111),
      .k9(32'b10111101100100101000011110001110)
  ) CON2D_118(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111000101011001011100101),
      .k2(32'b10111101101011000110110000101010),
      .k3(32'b10111100101010001100010111000111),
      .k4(32'b10111101100100101000010111011011),
      .k5(32'b10111101000100011111100001110011),
      .k6(32'b00111100000101110001010111010010),
      .k7(32'b10111101100110000011010011101110),
      .k8(32'b00111101111001011001111101111000),
      .k9(32'b10111100101011011110011000000011)
  ) CON2D_119(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010001100011010000011010),
      .k2(32'b00111101110000000001101101011000),
      .k3(32'b10111101111101101111011101010001),
      .k4(32'b00111101111000100011100100101000),
      .k5(32'b00111101101101101110010010010001),
      .k6(32'b10111100100000010100110100110011),
      .k7(32'b10111101101011011011000111100010),
      .k8(32'b00111100011001001001101001001010),
      .k9(32'b10111100001010010100111010111001)
  ) CON2D_120(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110011101111101110111110),
      .k2(32'b00111101110001011111100000111010),
      .k3(32'b10111101011111001001101100001101),
      .k4(32'b10111101111000011011110101101101),
      .k5(32'b00111101100001111110001011010100),
      .k6(32'b00111101000011010010001111100000),
      .k7(32'b10111101001100111010000010110011),
      .k8(32'b00111011000101110010000101111111),
      .k9(32'b10111101110010011111110110010011)
  ) CON2D_121(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100001001010101011100000110),
      .k2(32'b10111101110111101011110101110011),
      .k3(32'b10111100101000010000011011111110),
      .k4(32'b10111101110100011110110111011110),
      .k5(32'b10111101110011000011001000010010),
      .k6(32'b00111101110011010000110101111111),
      .k7(32'b00111101011100001110000001101100),
      .k8(32'b00111101011011001000110001100011),
      .k9(32'b00111100001110100100110010100000)
  ) CON2D_122(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011100010011011100000001101),
      .k2(32'b10111100100010001110010001010000),
      .k3(32'b10111101100001001111110101001010),
      .k4(32'b00111100110011010101111111100010),
      .k5(32'b10111100110001010010110010000101),
      .k6(32'b10111101101110101100001111011101),
      .k7(32'b10111100110111010001101111001010),
      .k8(32'b10111101011000101101111110001100),
      .k9(32'b10111011111010100111111001011001)
  ) CON2D_123(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000011111100110000010001),
      .k2(32'b10111100110000010111001000100111),
      .k3(32'b10111101001100010100011100000000),
      .k4(32'b10111101100100011110000001011100),
      .k5(32'b10111101101111110100010000110000),
      .k6(32'b00111101110010110001001011100001),
      .k7(32'b10111101001001000110010110111100),
      .k8(32'b00111100001000101110110011110011),
      .k9(32'b10111101101110101000010110110100)
  ) CON2D_124(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100100111011111001110100),
      .k2(32'b00111101010111111011101010000001),
      .k3(32'b00111101001011000011101001010001),
      .k4(32'b00111100101000000100010011111111),
      .k5(32'b00111101111001111100010110110011),
      .k6(32'b00111100011011001010101011100100),
      .k7(32'b10111101010110100010000111000110),
      .k8(32'b10111101001000110011111011000110),
      .k9(32'b10111011010111110110010100000000)
  ) CON2D_125(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100101010000010001010100),
      .k2(32'b00111100101011000110101111000111),
      .k3(32'b10111101111110011111111001000101),
      .k4(32'b10111101001011110100110110100000),
      .k5(32'b00111011101001100010110111101011),
      .k6(32'b10111101100101100110000001011000),
      .k7(32'b00111100101110100101010011111011),
      .k8(32'b10111101101010001111000101111100),
      .k9(32'b00111101010011100111010100001111)
  ) CON2D_126(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100010000100111110000),
      .k2(32'b10111100111001110100011011010011),
      .k3(32'b10111011110100000110111110100111),
      .k4(32'b00111101110011111001011110010100),
      .k5(32'b10111101100100010110010100010100),
      .k6(32'b10111100110000001001111001110111),
      .k7(32'b10111110000001110000011010000111),
      .k8(32'b00111101100000101111001011111110),
      .k9(32'b00111100011000011100010100110011)
  ) CON2D_127(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101001010011100100110001),
      .k2(32'b00111100110000011100100010001011),
      .k3(32'b10111101100011100111011011000100),
      .k4(32'b10111101110011100111011100101111),
      .k5(32'b00111101010101100001011100001100),
      .k6(32'b00111101101001001110110110010001),
      .k7(32'b10111101100101101000001001001100),
      .k8(32'b00111101000000010100100010110110),
      .k9(32'b00111100101101110111100001011001)
  ) CON2D_128(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[7][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111001000001000101000111110100)
)   op8(
    .i_pipeline_layer4(i_CORE_IP1[7]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*8-1:DATA_WIDTH*7])
);

/// CON2D_9///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111011100101101111111011),
      .k2(32'b00111101011100111100111101011100),
      .k3(32'b10111100111110111101010110011111),
      .k4(32'b00111101101111001000100010100111),
      .k5(32'b10111101001001100100010010001110),
      .k6(32'b10111101101101100011000010111100),
      .k7(32'b10111101011101100111010111101000),
      .k8(32'b00111101001011000001101011011011),
      .k9(32'b10111101100110011111000100001010)
  ) CON2D_129(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111010100000111011100000010000),
      .k2(32'b00111011100111110000110010110110),
      .k3(32'b00111101010111110011100100111111),
      .k4(32'b10111101000000011001100000001110),
      .k5(32'b10111101010101100101110100010001),
      .k6(32'b00111101110110010010110001000011),
      .k7(32'b00111101110001011011111101010110),
      .k8(32'b10111101101101110001011101000011),
      .k9(32'b00111101111111100001001000001110)
  ) CON2D_130(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110100101010000101010101),
      .k2(32'b10111100111011011100101001100001),
      .k3(32'b10111100011011011000111101000010),
      .k4(32'b00111101010110010011110001111111),
      .k5(32'b10111101001010001111010111100001),
      .k6(32'b00111101101011110110101110110100),
      .k7(32'b00111101100110110011011010101111),
      .k8(32'b10111101011110110010110100110110),
      .k9(32'b10111101110100001111011101010111)
  ) CON2D_131(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011101110000010100110000),
      .k2(32'b00111101001100010011111011010010),
      .k3(32'b00111101011000000001000001001010),
      .k4(32'b10111101100011010000000011110111),
      .k5(32'b00111101001011011001100011000000),
      .k6(32'b10111101101010010100000001011100),
      .k7(32'b10111001111111101001101100110000),
      .k8(32'b00111101100110001110000110101001),
      .k9(32'b10111100011001110100001100010101)
  ) CON2D_132(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000101001110001010001110),
      .k2(32'b00111101100101101010001101010111),
      .k3(32'b10111100001000011000100010111101),
      .k4(32'b10111101010101101101011011110110),
      .k5(32'b00111101110100100000111011011011),
      .k6(32'b00111101100010000111011101011110),
      .k7(32'b00111101001010011001101100010011),
      .k8(32'b10111101100010000000111110111100),
      .k9(32'b10111101100010011011111011101101)
  ) CON2D_133(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100001100010110010111100),
      .k2(32'b10111101101110101010100000000010),
      .k3(32'b10111101101010011110011011011111),
      .k4(32'b10111101100100010101110100100010),
      .k5(32'b10111101110100111010011001100100),
      .k6(32'b10111101010010000111111111110011),
      .k7(32'b00111100000101001111001011011000),
      .k8(32'b00111101000011010000000010000011),
      .k9(32'b00111101010111100010011010011001)
  ) CON2D_134(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101101001001101100101101),
      .k2(32'b10111101111100111010110101100001),
      .k3(32'b00111100011101100001100001110001),
      .k4(32'b10111101000001001010100101110100),
      .k5(32'b10111101100011101110111011010001),
      .k6(32'b00111101111000110001000110100010),
      .k7(32'b10111100010011000001101010110111),
      .k8(32'b00111101101101011110110001011000),
      .k9(32'b00111101110111000010000101010001)
  ) CON2D_135(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011100101111100011100010),
      .k2(32'b00111101010101111011010010100010),
      .k3(32'b10111101000111100010101000110101),
      .k4(32'b00111101101001100111010111001001),
      .k5(32'b10111100101001101000100111010100),
      .k6(32'b10111101100100101110011001111011),
      .k7(32'b10111101110011101100111101010100),
      .k8(32'b10111101010001111011001000111010),
      .k9(32'b10111100101101001001001000110110)
  ) CON2D_136(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110101001011110011010000),
      .k2(32'b00111101110011010110100011011100),
      .k3(32'b10111101100000001010101110000000),
      .k4(32'b10111101000110011010000110101011),
      .k5(32'b00111011110001111110000101101001),
      .k6(32'b10111101010000101011101101010001),
      .k7(32'b10111101001010010100010101110101),
      .k8(32'b10111101101001001110000100000001),
      .k9(32'b10111100111010011011100111010001)
  ) CON2D_137(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100111011010001101000100),
      .k2(32'b10111100100011110011101101101100),
      .k3(32'b00111101101011100001000100000000),
      .k4(32'b00111100000011001110101100111101),
      .k5(32'b00111101111011100111100101011011),
      .k6(32'b10111101101000101001000001101001),
      .k7(32'b00111100100110001110101111111001),
      .k8(32'b10111101110011100011000110001110),
      .k9(32'b10111101100000110110101000010011)
  ) CON2D_138(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010101011011011111110100),
      .k2(32'b10111100111000100110000000111111),
      .k3(32'b00111011101100010111001001111001),
      .k4(32'b00111101000100101101110001100001),
      .k5(32'b10111101101111101111000001010001),
      .k6(32'b10111101010100101011110110011010),
      .k7(32'b00111101100100101110110011010010),
      .k8(32'b00111101000011010010100100000000),
      .k9(32'b10111101110101000111100001000001)
  ) CON2D_139(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100100110011011000001101),
      .k2(32'b00111011111101101111001111101100),
      .k3(32'b00111101111100111000111000101000),
      .k4(32'b10111100111011111011110011110001),
      .k5(32'b00111101100001010101010000110100),
      .k6(32'b00111100110000000011110101111001),
      .k7(32'b00111101110001101011101110101100),
      .k8(32'b10111101100001000010000000111110),
      .k9(32'b00111101100011100101110100111101)
  ) CON2D_140(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001101001100110011101011),
      .k2(32'b10111101101100011011101011001001),
      .k3(32'b10111101111011101001110011001100),
      .k4(32'b10111011001110011101101000000010),
      .k5(32'b10111101101100111111100110101000),
      .k6(32'b00111011110101101000011101111101),
      .k7(32'b00111101111011001111011010101100),
      .k8(32'b10111100011000101011000110100001),
      .k9(32'b00111101111011111011100100100010)
  ) CON2D_141(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111110000001110011111100111100),
      .k2(32'b10111101111110100000011111010101),
      .k3(32'b00111011110010001101001111010101),
      .k4(32'b10111101010100100111010110011110),
      .k5(32'b00111011111110010010011111000001),
      .k6(32'b10111101110000110011000000101110),
      .k7(32'b10111110000011011110110001111111),
      .k8(32'b10111101001010110010101000010001),
      .k9(32'b10111101101010001111010111111111)
  ) CON2D_142(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011001110011110001000100),
      .k2(32'b10111101000111110010011101101000),
      .k3(32'b00111100011111110000001001000001),
      .k4(32'b00111101100110000111110101111110),
      .k5(32'b00111101011100000011111001001101),
      .k6(32'b10111101100011111010000110100101),
      .k7(32'b10111011011101101111110100000001),
      .k8(32'b00111101000000011110000011010001),
      .k9(32'b00111110000000011111000110110011)
  ) CON2D_143(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111000111000111101000110),
      .k2(32'b00111100001001111101100011111000),
      .k3(32'b10111101101100001101001100101001),
      .k4(32'b10111101110101110001101111000011),
      .k5(32'b00111100111000100111001011000111),
      .k6(32'b00111100100100001001110100110110),
      .k7(32'b10111110000000111111101111111101),
      .k8(32'b00111100001100011101101011111111),
      .k9(32'b10111101100001010110011010011100)
  ) CON2D_144(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[8][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100001011110110110011111010)
)   op9(
    .i_pipeline_layer4(i_CORE_IP1[8]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*9-1:DATA_WIDTH*8])
);

/// CON2D_10///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101010110001001000100010),
      .k2(32'b00111101010101011110110001000001),
      .k3(32'b00111101101111011101001011010010),
      .k4(32'b00111101001000010111011001001010),
      .k5(32'b00111101110110111010000111101011),
      .k6(32'b00111100100100100111101000110101),
      .k7(32'b00111101111001011111100000111100),
      .k8(32'b10111010101110010110001100100101),
      .k9(32'b00111101010111101001111000011011)
  ) CON2D_145(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101101011010101111001100),
      .k2(32'b10111101100000001010000110100011),
      .k3(32'b00111101000110110000001110000000),
      .k4(32'b10111101101000101000000101011100),
      .k5(32'b00111101011100001100010010101101),
      .k6(32'b10111101100011000110000010101000),
      .k7(32'b10111101010111110000111101000101),
      .k8(32'b00111101101101100100001000111100),
      .k9(32'b00111101110011010010010101000101)
  ) CON2D_146(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110001111101001000010010),
      .k2(32'b00111101100010110011110110010001),
      .k3(32'b00111100101010010110101111110010),
      .k4(32'b10111100100001010110100010010110),
      .k5(32'b10111101110101001111101100011000),
      .k6(32'b00111101000101101100000110010110),
      .k7(32'b10111011111111101000000001000001),
      .k8(32'b10111101100101111101001010010010),
      .k9(32'b10111101101101010100001110010101)
  ) CON2D_147(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110011100011100100101000),
      .k2(32'b00111100111111010111001111110000),
      .k3(32'b10111101011011100110001010010101),
      .k4(32'b10111101010001101001000101100000),
      .k5(32'b00111101101101011010110010111100),
      .k6(32'b10111100000111101000111110001011),
      .k7(32'b00111101101111111100110111111100),
      .k8(32'b10111101100000101111010000000000),
      .k9(32'b00111101011011101010010110001110)
  ) CON2D_148(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110101110011110011111001),
      .k2(32'b00111101101111101100110011101100),
      .k3(32'b10111101110111101110101011101011),
      .k4(32'b00111100010000110010000000000110),
      .k5(32'b10111100111110110001110000110001),
      .k6(32'b10111101101010101010000001100010),
      .k7(32'b10111101110000111010101100010110),
      .k8(32'b10111100101011101111011001110000),
      .k9(32'b10111101111100011101101110010111)
  ) CON2D_149(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111001010001001001100),
      .k2(32'b00111011100010101011000010001101),
      .k3(32'b10111101100010101110010001010100),
      .k4(32'b10111011110101100001010111000001),
      .k5(32'b00111101001001111111011011111110),
      .k6(32'b00111011111000010011000101011100),
      .k7(32'b10111100101010110011110011010010),
      .k8(32'b00111101011101101111000010100011),
      .k9(32'b10111101011001001110001111011010)
  ) CON2D_150(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001101111010011101001000),
      .k2(32'b00111101101101110010111000101010),
      .k3(32'b10111100010111111110001100011110),
      .k4(32'b10111101011100101011000001010010),
      .k5(32'b00111100100101110000000111010100),
      .k6(32'b10111101111110001110011111101101),
      .k7(32'b10111101001101100101001110000001),
      .k8(32'b10111101010110110110100110101101),
      .k9(32'b00111011111111001101101101110101)
  ) CON2D_151(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100001111111011000000111),
      .k2(32'b00111100110101101000011101011000),
      .k3(32'b10111100100010000110101111010000),
      .k4(32'b00111101010101100001101011101111),
      .k5(32'b00111101110100010110111010011011),
      .k6(32'b00111101110011110110110111010100),
      .k7(32'b00111101000111111010110000110100),
      .k8(32'b00111100010100010101011100011101),
      .k9(32'b10111010110011001110010110110011)
  ) CON2D_152(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110010000100100000110001),
      .k2(32'b10111101000010000001101100010100),
      .k3(32'b10111101110110000100111011110111),
      .k4(32'b10111101110011010001001000111000),
      .k5(32'b10111100011001011110011011001011),
      .k6(32'b10111101111110010000100100001000),
      .k7(32'b10111101001111100100110000000000),
      .k8(32'b00111101010011111100011000111001),
      .k9(32'b00111101110101011011101010000011)
  ) CON2D_153(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010010110011011001001000),
      .k2(32'b10111100100111000110111111011111),
      .k3(32'b00111100101100111000111100101101),
      .k4(32'b00111101001100001011100001000100),
      .k5(32'b10111100100100011001010001000010),
      .k6(32'b00111100001100001001111110100111),
      .k7(32'b00111101000010000011001010101000),
      .k8(32'b00111101101100111000010011010110),
      .k9(32'b10111101001001111100000010001100)
  ) CON2D_154(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001001001001000001011),
      .k2(32'b10111101010000110000011111000100),
      .k3(32'b10111101101101010110000000000101),
      .k4(32'b10111101110000111111110000101001),
      .k5(32'b10111101111010100011101100110100),
      .k6(32'b00111100111001101110000100100101),
      .k7(32'b10111100111011011010001011111011),
      .k8(32'b00111101010000001111001010111001),
      .k9(32'b00111101111001011010110100000100)
  ) CON2D_155(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100111011100000101110),
      .k2(32'b10111101101001110011000000001101),
      .k3(32'b10111101100001111111011000001010),
      .k4(32'b10111100011100001000100010010001),
      .k5(32'b10111101110101110011011100101101),
      .k6(32'b00111101110100100001000101101010),
      .k7(32'b10111101110011001100110111011111),
      .k8(32'b10111100010110111110000011011101),
      .k9(32'b10111101000111001010000101110101)
  ) CON2D_156(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111001001100101100011111),
      .k2(32'b10111010100110000000000011110001),
      .k3(32'b00111101101100001010111111100110),
      .k4(32'b00111101001100101000110000100110),
      .k5(32'b00111101100011010010001001010000),
      .k6(32'b00111101110011011010000111100011),
      .k7(32'b10111101110001100101000011111101),
      .k8(32'b10111101111011110110111111101110),
      .k9(32'b10111101100001011101110100111010)
  ) CON2D_157(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010001111111101101110101),
      .k2(32'b10111101000111110000111001101000),
      .k3(32'b00111100001111010001110111000011),
      .k4(32'b00111101000010110010101001100000),
      .k5(32'b00111101110010101100010011000000),
      .k6(32'b10111101101101111010101100111010),
      .k7(32'b00111101011101101100111100100110),
      .k8(32'b10111101110100001100001000011000),
      .k9(32'b10111100111000000011011100111011)
  ) CON2D_158(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101110001000011000001001),
      .k2(32'b10111101010010111010110101101000),
      .k3(32'b00111101111001011001001010010100),
      .k4(32'b10111101100011001000111011110101),
      .k5(32'b00111101111001111111000101101001),
      .k6(32'b10111101110011001111110100110100),
      .k7(32'b00111101110111101101011100100010),
      .k8(32'b00111101010010111010011110100111),
      .k9(32'b00111101101011100110010111000100)
  ) CON2D_159(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100000100110111000111),
      .k2(32'b10111100000010100101100011111010),
      .k3(32'b10111101011000001000000000100011),
      .k4(32'b00111101100011100100010010100000),
      .k5(32'b00111101100100010100000000111000),
      .k6(32'b10111101001000001000010111111101),
      .k7(32'b00111101110011100010110111011001),
      .k8(32'b00111100000110101110001001010100),
      .k9(32'b10111101101000010010001010011001)
  ) CON2D_160(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[9][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011111111001111011000000001)
)   op10(
    .i_pipeline_layer4(i_CORE_IP1[9]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*10-1:DATA_WIDTH*9])
);

/// CON2D_11///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100011110100110101111100),
      .k2(32'b00111101101000011111001100000110),
      .k3(32'b10111100110101111111010011010100),
      .k4(32'b10111100010001111001111111010101),
      .k5(32'b00111101100010101100001011000010),
      .k6(32'b00111101111011111101011100011000),
      .k7(32'b00111011111010111100110000001001),
      .k8(32'b10111101101100000110000111000011),
      .k9(32'b00111101001001100011100011001100)
  ) CON2D_161(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100001001110011001010011),
      .k2(32'b00111100111101011011111010001110),
      .k3(32'b00111101010111100111011110111001),
      .k4(32'b00111110000011010110000111001000),
      .k5(32'b10111100100111111000011010110011),
      .k6(32'b10111011001000001100000100011001),
      .k7(32'b00111101110100010011101011000001),
      .k8(32'b10111101110010101101010100010000),
      .k9(32'b10111101010101000110110001111101)
  ) CON2D_162(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100011110100001101011000),
      .k2(32'b00111101100011100100001100111001),
      .k3(32'b00111101110000010111111100001000),
      .k4(32'b10111100111000000000100111011001),
      .k5(32'b10111101101111110111000100010001),
      .k6(32'b00111101001001101110101101001111),
      .k7(32'b00111101110000111000010100001110),
      .k8(32'b00111101001000001100010111111101),
      .k9(32'b10111100010110100101111110010001)
  ) CON2D_163(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110011100110101000000100),
      .k2(32'b00111100001010101001100001111011),
      .k3(32'b10111101110111111111101100111001),
      .k4(32'b10111100100110010111100011100001),
      .k5(32'b10111101100100101111010111000000),
      .k6(32'b10111101001011011111011100101111),
      .k7(32'b10111100001011100100000000001010),
      .k8(32'b00111100100111011010001001001011),
      .k9(32'b10111101011001011001001000010000)
  ) CON2D_164(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100110101010011101001000),
      .k2(32'b00111101111011100110000011100011),
      .k3(32'b10111101011101110101111010000101),
      .k4(32'b10111101100001001010010101110010),
      .k5(32'b00111100010000011011111011010101),
      .k6(32'b00111110000000000011011111101101),
      .k7(32'b00111101011001110110100010110011),
      .k8(32'b00111101011101101111111101011111),
      .k9(32'b00111101100001001000001000110100)
  ) CON2D_165(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110000001011100101100111),
      .k2(32'b10111100011001101100101011010111),
      .k3(32'b10111100101111111110100011100101),
      .k4(32'b00111101110111100110000101011001),
      .k5(32'b00111101111010101000111001011111),
      .k6(32'b10111101101101000011010000101111),
      .k7(32'b00111100110101001001011100100000),
      .k8(32'b10111100111110111110010110011110),
      .k9(32'b10111101010001010010000111100111)
  ) CON2D_166(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111100101010000111111011),
      .k2(32'b10111101101111111111011011010001),
      .k3(32'b10111101000010100101110101111100),
      .k4(32'b00111101010000101101000010101011),
      .k5(32'b00111011011010101000110000011001),
      .k6(32'b00111101101000110010011100101011),
      .k7(32'b00111101100001011101100000101001),
      .k8(32'b10111011111011111101111101000000),
      .k9(32'b00111101010001101000011111101110)
  ) CON2D_167(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100110010100011110011111),
      .k2(32'b10111101100110010110011110100000),
      .k3(32'b00111100011100111001000000100111),
      .k4(32'b00111100101001001100010111111110),
      .k5(32'b10111101110000000000001101000001),
      .k6(32'b10111101101011111111111101010101),
      .k7(32'b10111101000101101100011001100001),
      .k8(32'b00111101000100000101010000111111),
      .k9(32'b10111101111001010001111000101010)
  ) CON2D_168(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100101011101111011111100),
      .k2(32'b10111101101011011101101011001100),
      .k3(32'b10111101011011011111010101010110),
      .k4(32'b10111011101111010100011111000111),
      .k5(32'b00111101110010000000001100010010),
      .k6(32'b00111101011011010010011110101000),
      .k7(32'b00111101111100110110000001001011),
      .k8(32'b10111101101101011111101101001111),
      .k9(32'b00111101001100110000110110010000)
  ) CON2D_169(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111101001010000000011111),
      .k2(32'b00111100001111100101100000000010),
      .k3(32'b00111101101001110010010001011101),
      .k4(32'b00111101110111001100001010101000),
      .k5(32'b00111101011101000001001011101101),
      .k6(32'b00111100100000011010111111000101),
      .k7(32'b00111101011101101110100100111100),
      .k8(32'b00111101110001100001010100001011),
      .k9(32'b00111101101111001001011100101010)
  ) CON2D_170(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110100010011011100110),
      .k2(32'b00111101011101111111010000101010),
      .k3(32'b00111101010100000001010011110100),
      .k4(32'b00111101110001101000111100111111),
      .k5(32'b00111011101010101010010110101110),
      .k6(32'b00111101001110011011100001000010),
      .k7(32'b00111010011110011010000100111000),
      .k8(32'b10111100101000100111001111100000),
      .k9(32'b10111101100001111100111010000101)
  ) CON2D_171(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100111011000101001001110),
      .k2(32'b00111101010110001011101010010001),
      .k3(32'b00111011101100101011111010111101),
      .k4(32'b00111101110001001001000011100101),
      .k5(32'b10111100111100010101101101010010),
      .k6(32'b00111101101001001110110101011110),
      .k7(32'b10111101000001110100001010011000),
      .k8(32'b00111101110110010010111101111101),
      .k9(32'b00111100100000100101101010100011)
  ) CON2D_172(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101010000101001100001100),
      .k2(32'b10111101110101010011001110011011),
      .k3(32'b10111101101001011111011010000101),
      .k4(32'b00111101000010101000110101101111),
      .k5(32'b10111101101000010001011001010100),
      .k6(32'b10111011101001100010100000111111),
      .k7(32'b10111011111101111010000110101000),
      .k8(32'b00111101001011111000011111111010),
      .k9(32'b10111101000011011011010011011001)
  ) CON2D_173(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000010010100100000010111),
      .k2(32'b00111101100101101101100100100011),
      .k3(32'b10111100111010110100010010100110),
      .k4(32'b00111011100011011011101010011001),
      .k5(32'b10111101110010101110111110110000),
      .k6(32'b00111101010001111010110111000110),
      .k7(32'b10111101011110010111010101111010),
      .k8(32'b10111101111100001111100010001010),
      .k9(32'b00111101000010000111111000000100)
  ) CON2D_174(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101010110000000100110100),
      .k2(32'b10111101101001100111000000010000),
      .k3(32'b10111110000001110011111100101100),
      .k4(32'b10111100110011101000111101101111),
      .k5(32'b00111101101110010011011011000111),
      .k6(32'b00111101001100001010110000000100),
      .k7(32'b10111101001011101000001101000000),
      .k8(32'b10111101010111010111010000101000),
      .k9(32'b10111110000000111001001011110111)
  ) CON2D_175(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100100100010000000110101),
      .k2(32'b10111101110000001111001000010100),
      .k3(32'b10111101010101000101110001101011),
      .k4(32'b10111100100111011011101010011110),
      .k5(32'b00111101101110011000010101100000),
      .k6(32'b00111101001001001001111010001011),
      .k7(32'b00111101000010110011000101000110),
      .k8(32'b10111100100000000111001010111110),
      .k9(32'b10111101001011101100001110111000)
  ) CON2D_176(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[10][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011101101111001110110111001)
)   op11(
    .i_pipeline_layer4(i_CORE_IP1[10]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*11-1:DATA_WIDTH*10])
);

/// CON2D_12///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001000011010100010100100),
      .k2(32'b00111100110001111101011011101110),
      .k3(32'b10111101001010111111100001110000),
      .k4(32'b10111101101110001011001100111000),
      .k5(32'b00111100101111110110011111100101),
      .k6(32'b00111100100011001101000001000011),
      .k7(32'b10111011101010001010110100110010),
      .k8(32'b10111101110111000000010010110001),
      .k9(32'b00111101111000011011000101010000)
  ) CON2D_177(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010001101011010001110001),
      .k2(32'b00111101011100101100101100000000),
      .k3(32'b10111101110001001111100101011001),
      .k4(32'b10111101011111000110111011011011),
      .k5(32'b00111101011001010010101001100101),
      .k6(32'b10111100101101100101101111100100),
      .k7(32'b10111011101111111000110111011011),
      .k8(32'b10111101111000000110011101010111),
      .k9(32'b10111101001101100001011001011101)
  ) CON2D_178(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011101100101000101000100100),
      .k2(32'b00111101101010000001100001111000),
      .k3(32'b10111101101011001100111001101010),
      .k4(32'b00111101100110011011010010000110),
      .k5(32'b10111100100100001011001111110111),
      .k6(32'b00111101000100111100110110001101),
      .k7(32'b00111101000110100011001101111110),
      .k8(32'b00111101001110110011101011111001),
      .k9(32'b10111101100110011000111100110110)
  ) CON2D_179(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111001011110001000000010101010),
      .k2(32'b10111101001110001110011001110000),
      .k3(32'b10111101101101011000000010110000),
      .k4(32'b10111100101100000111101011000111),
      .k5(32'b10111101101001010000011101100100),
      .k6(32'b00111101111011010011000101010111),
      .k7(32'b00111100111101110110101010101011),
      .k8(32'b10111101111011111101001000010111),
      .k9(32'b00111101110100100100000110011101)
  ) CON2D_180(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101110001111110101010000),
      .k2(32'b00111101101010000110111101001110),
      .k3(32'b00111011001001110101011011111101),
      .k4(32'b10111101101001010111110010100000),
      .k5(32'b10111100101011101101011100001111),
      .k6(32'b10111101111011001111011000011011),
      .k7(32'b00111011100011010010110111001100),
      .k8(32'b00111100101011100001010100011100),
      .k9(32'b00111101110101000110110101110100)
  ) CON2D_181(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101010011110111011111100),
      .k2(32'b10111101111000001010111100001110),
      .k3(32'b10111101001011010001011011000010),
      .k4(32'b10111101011010011000111011111011),
      .k5(32'b00111101100010010101000010001100),
      .k6(32'b00111011111100010110111100110111),
      .k7(32'b10111101001011001011011111011111),
      .k8(32'b10111100100110100100101101011110),
      .k9(32'b10111101101100110010010100101110)
  ) CON2D_182(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111110000011000010110010111101),
      .k2(32'b10111101101010101101111010110011),
      .k3(32'b00111101000111000011010010110111),
      .k4(32'b10111101110110001100110100000010),
      .k5(32'b00111101110001011000001101011000),
      .k6(32'b10111101101001111111000001101101),
      .k7(32'b10111101111100110111011111111000),
      .k8(32'b00111101110010010100010000011010),
      .k9(32'b10111101001001001110010000011111)
  ) CON2D_183(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100110010100110010100101101),
      .k2(32'b00111101111011010001101000111000),
      .k3(32'b10111101110110110111010010101111),
      .k4(32'b00111101111010100101111101110100),
      .k5(32'b00111101011010110011011110100111),
      .k6(32'b10111010100010011001011101100110),
      .k7(32'b00111101111100010101110110101000),
      .k8(32'b10111100100000010010001110101101),
      .k9(32'b10111100011001110100100010011101)
  ) CON2D_184(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100001000000010000101010),
      .k2(32'b10111101101011101110111111110100),
      .k3(32'b10111101011101111010100001000011),
      .k4(32'b00111100110111001000011011010000),
      .k5(32'b10111101110001100111111111001101),
      .k6(32'b10111101010001001111001100010101),
      .k7(32'b10111100111011011011111010100110),
      .k8(32'b10111100111110010101100001001111),
      .k9(32'b10111101100110001110111100101111)
  ) CON2D_185(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011100000111101010111000100),
      .k2(32'b00111100110111111001100011011111),
      .k3(32'b00111101110000100010100101111110),
      .k4(32'b10111101110011010101111001111110),
      .k5(32'b00111100101110001101010011000000),
      .k6(32'b00111101100100001111010110100001),
      .k7(32'b00111101111111001110110101000010),
      .k8(32'b00111101001000101100010101100111),
      .k9(32'b10111101110101001001101111100001)
  ) CON2D_186(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001011101010000000110),
      .k2(32'b10111101010011000101000010010100),
      .k3(32'b10111100110111100100100011011010),
      .k4(32'b10111101011100110010110111001010),
      .k5(32'b00111101100010010010110110001110),
      .k6(32'b00111101100111001010000101100010),
      .k7(32'b00111101110000010110000110111001),
      .k8(32'b10111011111101110011001001110010),
      .k9(32'b00111101001000010100011010101110)
  ) CON2D_187(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101111001000011001011101),
      .k2(32'b10111011011101001010001010111110),
      .k3(32'b10111101111101000001011010010000),
      .k4(32'b10111101011110010001100010101100),
      .k5(32'b10111101101001101000110011101110),
      .k6(32'b00111101010010011001111101000001),
      .k7(32'b10111100111101111001000101001101),
      .k8(32'b00111101101110010011111101100100),
      .k9(32'b10111101010001100101000011011111)
  ) CON2D_188(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011111111000101000100000010),
      .k2(32'b00111101101001011011101110111111),
      .k3(32'b10111101100100001110010100000101),
      .k4(32'b10111101111000011000101001001011),
      .k5(32'b10111101101000110111111111010001),
      .k6(32'b00111100111010000101101101111101),
      .k7(32'b00111100011111111110101011101001),
      .k8(32'b00111101001111110111111101001101),
      .k9(32'b00111101100101111101110001110111)
  ) CON2D_189(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111010001010111100001111),
      .k2(32'b00111100101101001010001100010110),
      .k3(32'b00111101000100111111100101101000),
      .k4(32'b10111100101111001011010111111101),
      .k5(32'b00111101000100110000011110000011),
      .k6(32'b10111101011001001001110101100100),
      .k7(32'b00111101011100001000011101010110),
      .k8(32'b10111101011001110011001000010001),
      .k9(32'b10111101000111110010101100100101)
  ) CON2D_190(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001000100101111100111),
      .k2(32'b00111101100110101100111111101000),
      .k3(32'b10111101110010111110000000011000),
      .k4(32'b10111100100111111000100011100111),
      .k5(32'b00111100010110101011101000011110),
      .k6(32'b00111101110000110110010011100101),
      .k7(32'b00111100101100101010101011001110),
      .k8(32'b00111100111100110100101100011010),
      .k9(32'b10111101101001011000010111010011)
  ) CON2D_191(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111101001100110110001101),
      .k2(32'b00111101110110010011010011100100),
      .k3(32'b10111101001111010000100010111110),
      .k4(32'b00111100111001011010001111001100),
      .k5(32'b00111101111000000111001011000000),
      .k6(32'b10111101100000101011000001000001),
      .k7(32'b00111100101000100100001100110111),
      .k8(32'b00111011010010111110000011111100),
      .k9(32'b00111101000011001111101001011010)
  ) CON2D_192(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[11][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111010001001010111011100111111)
)   op12(
    .i_pipeline_layer4(i_CORE_IP1[11]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*12-1:DATA_WIDTH*11])
);

/// CON2D_13///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011011100110101110100100111),
      .k2(32'b00111101101000010100000011111111),
      .k3(32'b10111100011010000010011011111000),
      .k4(32'b00111101010100101110101000100010),
      .k5(32'b10111011000110000100010101001101),
      .k6(32'b00111101001010000100001011100111),
      .k7(32'b00111100100011011010110110001100),
      .k8(32'b10111101001110010100001100011111),
      .k9(32'b00111100100000111100111101011001)
  ) CON2D_193(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110110111111000111111111),
      .k2(32'b10111101011111100100110111001111),
      .k3(32'b00111101100111100110101101110101),
      .k4(32'b10111101000011111100111101010010),
      .k5(32'b10111100011101001010000000111110),
      .k6(32'b10111101010000000100010010001011),
      .k7(32'b10111101101010111110001100011010),
      .k8(32'b00111101110010010001010000011110),
      .k9(32'b10111101011111111110001001101001)
  ) CON2D_194(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000010011110100110000011),
      .k2(32'b10111101110001110011011011101100),
      .k3(32'b00111101110110111000011100110100),
      .k4(32'b10111101001001000010001111100100),
      .k5(32'b10111101110100110010110001001110),
      .k6(32'b10111100111010100101011010110100),
      .k7(32'b00111101110001111101101100001101),
      .k8(32'b10111100101011100101110101011000),
      .k9(32'b00111101001000000110010010010111)
  ) CON2D_195(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100001011101001110011111001),
      .k2(32'b00111101110110010100101011100011),
      .k3(32'b00111101100001011100100100010110),
      .k4(32'b10111101111100011000001010001111),
      .k5(32'b10111101101011001001010000011101),
      .k6(32'b10111001100101001001110111110001),
      .k7(32'b10111101111001010111111000110101),
      .k8(32'b10111101111001100000010011010100),
      .k9(32'b00111100110011000111000110000111)
  ) CON2D_196(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100101000100101001100010),
      .k2(32'b10111101001000011111010001000100),
      .k3(32'b00111101101100010110101110011101),
      .k4(32'b00111101110110010111101110110100),
      .k5(32'b10111101101001100000001000000111),
      .k6(32'b00111101100010100110010001110010),
      .k7(32'b00111101001111100001101011001101),
      .k8(32'b10111101101110010011111001110101),
      .k9(32'b10111101101011100100111100101001)
  ) CON2D_197(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011110011011111101100001001),
      .k2(32'b00111100101010100011001000000100),
      .k3(32'b00111101000011011111001010110110),
      .k4(32'b00111101110111111011101001100010),
      .k5(32'b00111101100000111000111001001101),
      .k6(32'b00111101001110000000100100101011),
      .k7(32'b10111101100111101101111011011111),
      .k8(32'b00111100000100010100011011101100),
      .k9(32'b00111101000110001011110111101111)
  ) CON2D_198(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011101101100000000010000010),
      .k2(32'b00111110000000010101000110101111),
      .k3(32'b00111101110101011010100010111010),
      .k4(32'b00111110000000100011110110100111),
      .k5(32'b00111100011010000000011011010001),
      .k6(32'b00111101011000111100101101010110),
      .k7(32'b00111101100000110001111001001111),
      .k8(32'b00111101011000100111110000100111),
      .k9(32'b00111101011000100011101001011010)
  ) CON2D_199(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011111110111111010111011),
      .k2(32'b10111101010010110000010010110101),
      .k3(32'b00111101101010010101101011001100),
      .k4(32'b00111101101001101001000101101111),
      .k5(32'b10111101101111001100000010000110),
      .k6(32'b00111010111110111011111010101110),
      .k7(32'b00111101001000001111111110010011),
      .k8(32'b10111100111100110001111110010010),
      .k9(32'b00111101101111011011110111101110)
  ) CON2D_200(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110011101000001000111001),
      .k2(32'b10111100110010001100101011110101),
      .k3(32'b00111101111100111001100101101011),
      .k4(32'b00111101011000111111010000010000),
      .k5(32'b10111101110100011101110100010100),
      .k6(32'b10111101001110010010100000110010),
      .k7(32'b10111101110001001011001011011011),
      .k8(32'b00111100100110000011110011100001),
      .k9(32'b10111100101100111111101111000111)
  ) CON2D_201(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110101011100010011011010),
      .k2(32'b10111101111001001101001001101001),
      .k3(32'b00111101100000000010000110011010),
      .k4(32'b00111101100010010011110111111110),
      .k5(32'b00111101110101001111110010000111),
      .k6(32'b00111101110001000001110111111001),
      .k7(32'b10111101101010010011110110001011),
      .k8(32'b00111101100101011010000001111110),
      .k9(32'b10111101100101010011010110000111)
  ) CON2D_202(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010010110010111110101000),
      .k2(32'b10111101110100101111000011010111),
      .k3(32'b10111101111000101110110011111110),
      .k4(32'b00111101011001110010100110001010),
      .k5(32'b00111101111010000010001100110101),
      .k6(32'b00111101101000010000111111111011),
      .k7(32'b10111101000111000000100001001110),
      .k8(32'b00111101101011111011101000110110),
      .k9(32'b10111101110011000011001011100111)
  ) CON2D_203(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000001001110100011001100),
      .k2(32'b10111101110100011011000001110101),
      .k3(32'b10111101110100000000100111100010),
      .k4(32'b10111101011001111000111000011110),
      .k5(32'b00111011000000011011101001111101),
      .k6(32'b00111100100001101010011000011110),
      .k7(32'b00111101001100111101111001100001),
      .k8(32'b00111101101001010010110101110111),
      .k9(32'b00111100100110101010010101111100)
  ) CON2D_204(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011000100101100100000),
      .k2(32'b00111101011000100001110000001000),
      .k3(32'b00111101000100011010011010000000),
      .k4(32'b00111101110010010110100010101101),
      .k5(32'b00111100100101011001010101011110),
      .k6(32'b00111101101001001101011100001100),
      .k7(32'b10111100010001010011101111011100),
      .k8(32'b10111101010011011111000100011101),
      .k9(32'b00111101100101100001100011110010)
  ) CON2D_205(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011110011110101110011011010),
      .k2(32'b10111101111011100011001111011001),
      .k3(32'b00111101101110001000001100001101),
      .k4(32'b10111101110001100110010101010100),
      .k5(32'b00111100001001001100111110100001),
      .k6(32'b10111101110011011010110101111001),
      .k7(32'b00111101110001010001101101011101),
      .k8(32'b00111101111010101111100010111011),
      .k9(32'b10111101010101111011111100011011)
  ) CON2D_206(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100000011100001000101100110),
      .k2(32'b10111101110010011010001101010000),
      .k3(32'b00111100010100000000010001011110),
      .k4(32'b00111011110001101010110100001111),
      .k5(32'b10111101111101001000010010010001),
      .k6(32'b00111101011011010100000100110111),
      .k7(32'b10111101011110011100010001001111),
      .k8(32'b10111101100111011101011110110001),
      .k9(32'b10111101011110111101010101100000)
  ) CON2D_207(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100010101111100101011011111),
      .k2(32'b10111101100100111110011000000111),
      .k3(32'b10111101100110101111110110010011),
      .k4(32'b00111010111000101110011101100001),
      .k5(32'b00111101011000011011011100101100),
      .k6(32'b10111100111001011011001100011111),
      .k7(32'b10111101001010010100110101011011),
      .k8(32'b00111101111011000110110101100001),
      .k9(32'b00111101101111110111010110101100)
  ) CON2D_208(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[12][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011101000000111111110011011)
)   op13(
    .i_pipeline_layer4(i_CORE_IP1[12]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*13-1:DATA_WIDTH*12])
);

/// CON2D_14///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101001010011100101111001),
      .k2(32'b00111100010010011010001100110110),
      .k3(32'b00111101101001000010011101100101),
      .k4(32'b00111101101111111001110110100100),
      .k5(32'b10111101110011001110101011001001),
      .k6(32'b00111101111100101001111100000111),
      .k7(32'b10111101011110110101111111111111),
      .k8(32'b10111100111100111011110000011110),
      .k9(32'b10111101100101000111111000110111)
  ) CON2D_209(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001010000101100110100010),
      .k2(32'b10111101010110111010100011110101),
      .k3(32'b10111100110001010101011100000000),
      .k4(32'b10111101110010010110001100001010),
      .k5(32'b10111101101001111100001110101011),
      .k6(32'b00111101000110001101110111001101),
      .k7(32'b10111101001101011001110011100110),
      .k8(32'b10111011110100110010100100100110),
      .k9(32'b00111100100000011111101111001001)
  ) CON2D_210(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101010111000110001010001),
      .k2(32'b10111101110001111110001100100011),
      .k3(32'b00111101110111100110101001001110),
      .k4(32'b00111101100110110101000101100010),
      .k5(32'b10111101111001101000100101111000),
      .k6(32'b10111101010101000100110111000100),
      .k7(32'b10111101101000110110011000111011),
      .k8(32'b00111101110110011001001000100001),
      .k9(32'b00111101101101101010001000010101)
  ) CON2D_211(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101101100001001010010011),
      .k2(32'b10111101110110110001111011101000),
      .k3(32'b00111101110100110100011001100111),
      .k4(32'b10111100101011110110111001111111),
      .k5(32'b00111101110000011111000111101100),
      .k6(32'b00111101110110001110011000001000),
      .k7(32'b00111101110111001100100101111100),
      .k8(32'b10111100110100011100001010110011),
      .k9(32'b10111101110010110111000110011011)
  ) CON2D_212(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101000001111000110101011),
      .k2(32'b10111101110001011010111001011010),
      .k3(32'b00111100101101110010010110000111),
      .k4(32'b10111100101000101010010011010111),
      .k5(32'b00111101110101110100011010000100),
      .k6(32'b10111100100001110011101100010010),
      .k7(32'b10111101000101110110010001011111),
      .k8(32'b10111101111100001010101100001011),
      .k9(32'b00111101110100101110001100001101)
  ) CON2D_213(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111011000010101101001100),
      .k2(32'b00111101100000000011011100000000),
      .k3(32'b10111101101010100010000101101101),
      .k4(32'b10111101011001100001000110111100),
      .k5(32'b10111101011001111111110001000000),
      .k6(32'b10111101011000100111101000001111),
      .k7(32'b10111100111101100011110011100101),
      .k8(32'b10111101001001010001010101101000),
      .k9(32'b10111101100000000001011011000111)
  ) CON2D_214(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111100001010100011110),
      .k2(32'b10111101101100001110101111000101),
      .k3(32'b10111101110110100010111011011100),
      .k4(32'b00111101110010000011110001100101),
      .k5(32'b00111101110011011001010010110011),
      .k6(32'b00111100111000011111111011110101),
      .k7(32'b00111101010010001011000010111110),
      .k8(32'b00111011101000100100111101110011),
      .k9(32'b10111101000010010101111101100011)
  ) CON2D_215(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011111100100100101100111),
      .k2(32'b10111101110111001011111000100100),
      .k3(32'b00111101000101001001001100110101),
      .k4(32'b10111101010000011011111000000011),
      .k5(32'b10111100100001001101011011101011),
      .k6(32'b10111100010100100000001011011001),
      .k7(32'b00111101111100001111010111011001),
      .k8(32'b10111100011111011000101010001101),
      .k9(32'b10111101010010000101011111110011)
  ) CON2D_216(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110110000010010101010),
      .k2(32'b00111101000101111110111001001110),
      .k3(32'b10111101011011110101011011000110),
      .k4(32'b00111101011011100001000110111010),
      .k5(32'b00111101010110000111000010011001),
      .k6(32'b10111101001101000011011110001001),
      .k7(32'b10111101111110111111011110111100),
      .k8(32'b10111101000001010000100010011000),
      .k9(32'b10111100111100111111000010110001)
  ) CON2D_217(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111101110010001001100101),
      .k2(32'b10111011100011101111010110011000),
      .k3(32'b10111101101110011110111000101101),
      .k4(32'b00111101111100011000111001110010),
      .k5(32'b10111101101001000010100101011001),
      .k6(32'b10111100111111100001101001100111),
      .k7(32'b10111011100110100110000110011110),
      .k8(32'b00111101100000100001101011010000),
      .k9(32'b10111010011101001100000010011111)
  ) CON2D_218(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000011010110111011010010),
      .k2(32'b00111101010010111101111101001101),
      .k3(32'b00111101010000111010001011111001),
      .k4(32'b10111100110101100110001100110100),
      .k5(32'b10111101110010100001011001101110),
      .k6(32'b10111101100100001111101110010000),
      .k7(32'b00111101110111101001111111110011),
      .k8(32'b10111101111001010001011011101000),
      .k9(32'b10111101110111011001101010101000)
  ) CON2D_219(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111110011001001101110101),
      .k2(32'b10111101100100001000110100111101),
      .k3(32'b00111100100001010111101100100111),
      .k4(32'b10111101110010111001011100010010),
      .k5(32'b10111101111100111011000111101101),
      .k6(32'b10111101111110011000110111110101),
      .k7(32'b10111101100100110111111000000100),
      .k8(32'b10111101111110001000110100101111),
      .k9(32'b00111101011000011101011110110000)
  ) CON2D_220(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100110101010001111001010011),
      .k2(32'b00111100101100000011001100000110),
      .k3(32'b10111101010111000011111011111010),
      .k4(32'b00111101101000000111111110001111),
      .k5(32'b10111100100110100010100111001000),
      .k6(32'b00111101011100001100001000111000),
      .k7(32'b00111101101010010101101010011100),
      .k8(32'b00111101110101101110100010011100),
      .k9(32'b10111101101000011000000100101000)
  ) CON2D_221(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000111100010100010001101),
      .k2(32'b00111101111110100100111001110100),
      .k3(32'b10111011100010011110110000001000),
      .k4(32'b00111101100111110100111000110000),
      .k5(32'b00111101100010001010101010100011),
      .k6(32'b00111101100000010101000010001001),
      .k7(32'b10111101101011000110001011011010),
      .k8(32'b10111101101110101000110011101101),
      .k9(32'b00111101001000111010111010001111)
  ) CON2D_222(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011000000010101010001000101),
      .k2(32'b00111100100011110101011111011011),
      .k3(32'b10111101000011011110111110101000),
      .k4(32'b10111101010000100000010011001000),
      .k5(32'b00111100011110100001111011010110),
      .k6(32'b00111101110100001110010010101111),
      .k7(32'b00111100111110111000100010011010),
      .k8(32'b10111100101101011011010010100101),
      .k9(32'b00111101110100010111100110101111)
  ) CON2D_223(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110000100001100110100110),
      .k2(32'b00111101110011001100000011110000),
      .k3(32'b00111101110001101101111001101010),
      .k4(32'b10111011101100100100111000011100),
      .k5(32'b10111101010110010110010011101110),
      .k6(32'b10111101010110001101101000010001),
      .k7(32'b10111101100000110010111111101101),
      .k8(32'b00111100000011011010101110000000),
      .k9(32'b00111101111011011001010110011100)
  ) CON2D_224(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[13][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111010111001100011111001110101)
)   op14(
    .i_pipeline_layer4(i_CORE_IP1[13]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*14-1:DATA_WIDTH*13])
);

/// CON2D_15///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111101001000101001111100),
      .k2(32'b00111101000101000100111011110111),
      .k3(32'b00111011111010000101111100010111),
      .k4(32'b10111101010111011111110001001101),
      .k5(32'b00111101100110001000000001010011),
      .k6(32'b00111101101111001000110011000000),
      .k7(32'b10111101000111110100011011000001),
      .k8(32'b00111101111010010100100000000000),
      .k9(32'b00111100110110010011001010001011)
  ) CON2D_225(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011100001111010000000111),
      .k2(32'b10111100110011011110110111010110),
      .k3(32'b00111110000000111001111100100001),
      .k4(32'b10111011101011100100101101000010),
      .k5(32'b10111101100000100100110100011111),
      .k6(32'b00111110000100110001011101110010),
      .k7(32'b10111101010001000001110110110110),
      .k8(32'b00111101100101001111110111111011),
      .k9(32'b00111101110110101000001001100010)
  ) CON2D_226(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101010111111010011110011),
      .k2(32'b10111101100111001111111001100111),
      .k3(32'b10111101010111100100001010000100),
      .k4(32'b00111011111100101000100011101001),
      .k5(32'b10111101111101011000010110001011),
      .k6(32'b10111011101010110001100001000000),
      .k7(32'b00111011010001101111001001110001),
      .k8(32'b10111101101000001100001111011011),
      .k9(32'b10111101001011000000100001001001)
  ) CON2D_227(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000110110011101001111101),
      .k2(32'b10111101011101011110111110001000),
      .k3(32'b00111100110110010110010100110111),
      .k4(32'b10111101010100000101010100101101),
      .k5(32'b10111100100100010000110011001000),
      .k6(32'b10111101100000000000100001001111),
      .k7(32'b00111001100110001100101011000101),
      .k8(32'b10111101100010101101001001111010),
      .k9(32'b00111101110110101110001001010111)
  ) CON2D_228(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100000100100111010011100),
      .k2(32'b00111101001100111000000100100010),
      .k3(32'b10111101111011001100011101101010),
      .k4(32'b10111101110011111010101001101101),
      .k5(32'b10111101100001011001010001110011),
      .k6(32'b10111100100101100100011111001001),
      .k7(32'b00111100110001101000000000000110),
      .k8(32'b00111101011101000101110111100101),
      .k9(32'b10111101111000000100011101010010)
  ) CON2D_229(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110000111000111100111000),
      .k2(32'b00111100101011010111100111001110),
      .k3(32'b10111101101111111101101100001011),
      .k4(32'b10111101101111110010011111010110),
      .k5(32'b10111101111100111111110101011100),
      .k6(32'b00111100100100011010000111000010),
      .k7(32'b10111101111111001001101000100101),
      .k8(32'b10111101100011100001011000100000),
      .k9(32'b10111101100001101100111101111000)
  ) CON2D_230(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101010010000110010101001),
      .k2(32'b10111100100000100000101100000100),
      .k3(32'b10111101100100100011101101100011),
      .k4(32'b10111101100110010010101000111111),
      .k5(32'b10111101010001011111011011011100),
      .k6(32'b10111101001110011111010000111111),
      .k7(32'b10111101010011101011010111001100),
      .k8(32'b00111101100111001001111010010110),
      .k9(32'b10111101000111100001011110001001)
  ) CON2D_231(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100001100000001110000101011),
      .k2(32'b00111101100000011011000110011000),
      .k3(32'b00111101110111001100010011110000),
      .k4(32'b00111101110000101111110000010000),
      .k5(32'b10111101011000111010100000110010),
      .k6(32'b00111100101111000010111001000000),
      .k7(32'b00111100001010011010110110110010),
      .k8(32'b10111101000111010101010001001010),
      .k9(32'b00111101010101010001010100001100)
  ) CON2D_232(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011010010101011110110011),
      .k2(32'b10111101100011111111010000100111),
      .k3(32'b10111100100011111111010101000001),
      .k4(32'b00111101110010100011001000111001),
      .k5(32'b10111100010101101110101111011111),
      .k6(32'b10111010111100001001010100111111),
      .k7(32'b00111101101010111011111111100110),
      .k8(32'b00111101110001110111001111010101),
      .k9(32'b00111101101111101100001011000100)
  ) CON2D_233(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001011100001101011101),
      .k2(32'b00111101000000000110010001111001),
      .k3(32'b10111100100011100111110001000001),
      .k4(32'b10111101100010001101111011000101),
      .k5(32'b10111101101011100111111111100111),
      .k6(32'b10111101101111110100110110001101),
      .k7(32'b10111101000101100110111010100100),
      .k8(32'b00111101101101001101011111100101),
      .k9(32'b00111101110100011000111000101101)
  ) CON2D_234(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100010111001110011101111),
      .k2(32'b10111100010011111001011100011100),
      .k3(32'b00111101100000011011100111100001),
      .k4(32'b10111101101000001010010010010100),
      .k5(32'b00111101101010110110010111100111),
      .k6(32'b00111100001101101100011101100011),
      .k7(32'b10111101000110101111101010010111),
      .k8(32'b10111101000010000110000000110000),
      .k9(32'b10111101000000001000111101001101)
  ) CON2D_235(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100001000110000101000011011),
      .k2(32'b10111101010110001001001011011010),
      .k3(32'b00111101010001111110101000010111),
      .k4(32'b00111101101110100111110110101110),
      .k5(32'b10111101001110110110010111000110),
      .k6(32'b10111011001100100010010011000011),
      .k7(32'b10111101101110100001101111011011),
      .k8(32'b10111101000111001100011100100111),
      .k9(32'b00111101001001011110011111011111)
  ) CON2D_236(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011011011101011101111000),
      .k2(32'b10111100100011011001110101001001),
      .k3(32'b10111101100010000001011100000101),
      .k4(32'b10111101111001100100110000110011),
      .k5(32'b00111101100101110001011000010001),
      .k6(32'b10111101100001010110001011001000),
      .k7(32'b10111100100000110000100011000000),
      .k8(32'b10111101000110000100010100011000),
      .k9(32'b10111101101101110100110010110111)
  ) CON2D_237(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001110001001111101010011),
      .k2(32'b10111100100100101100001101101111),
      .k3(32'b00111100100110100000011011000010),
      .k4(32'b10111100001000011010110101100110),
      .k5(32'b00111101110100001010101000000100),
      .k6(32'b10111101100001111101111101111000),
      .k7(32'b00111010101011001000001010101001),
      .k8(32'b10111100111001001101111110001001),
      .k9(32'b10111101101010011100111111111101)
  ) CON2D_238(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111011100101010011110101),
      .k2(32'b00111101100100110110100010100100),
      .k3(32'b00111101110111110010010110111001),
      .k4(32'b00111100000011101100100100011101),
      .k5(32'b10111101100000100001011000000110),
      .k6(32'b00111101110111101011110110001100),
      .k7(32'b10111101100111000001100011000111),
      .k8(32'b10111101100001101111001010101001),
      .k9(32'b00111101010010000100100011010001)
  ) CON2D_239(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100010111011111100001100100),
      .k2(32'b10111011110010011111100111001101),
      .k3(32'b10111101111110011011110111001101),
      .k4(32'b10111101000110101011101000100011),
      .k5(32'b10111011100010010000111111000011),
      .k6(32'b00111101100100001000011010111000),
      .k7(32'b00111100000011110011001101111110),
      .k8(32'b00111101110000110010010110011111),
      .k9(32'b00111010001010001001010000101010)
  ) CON2D_240(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[14][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111001110011011111011010101111)
)   op15(
    .i_pipeline_layer4(i_CORE_IP1[14]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*15-1:DATA_WIDTH*14])
);

/// CON2D_16///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011110111111100001010111),
      .k2(32'b00111101110111011110100001100011),
      .k3(32'b10111100001011111111010111101001),
      .k4(32'b10111100100010111011111101001011),
      .k5(32'b10111101101001011101001011110000),
      .k6(32'b00111101110000111100011111001000),
      .k7(32'b00111100000110110100000010101101),
      .k8(32'b10111100110001111100101101010011),
      .k9(32'b10111101001110100001011000000101)
  ) CON2D_241(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011010010010110000100111),
      .k2(32'b00111101000011011001110001010111),
      .k3(32'b10111100111011011000010000011010),
      .k4(32'b10111101101101110011001011000100),
      .k5(32'b10111010111100110100001101000001),
      .k6(32'b00111100111111001010010101010000),
      .k7(32'b00111101110001011100101111000110),
      .k8(32'b00111101101111000100100011000010),
      .k9(32'b10111101001110101110111110001011)
  ) CON2D_242(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111000000010001110100000),
      .k2(32'b10111101100001110111100100101010),
      .k3(32'b10111101110101000110111110101010),
      .k4(32'b10111100010111110101011100110100),
      .k5(32'b00111101000101111101101101101011),
      .k6(32'b00111011111100001100010001010110),
      .k7(32'b10111101101010011001110000101000),
      .k8(32'b00111101001111110000011101000101),
      .k9(32'b00111011111101011001111001001011)
  ) CON2D_243(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111011000001011010111000),
      .k2(32'b00111101100111011111011101110001),
      .k3(32'b10111101101111011010001100000100),
      .k4(32'b00111101100001100011010101001111),
      .k5(32'b10111101001110010100011000000111),
      .k6(32'b00111100111111001101110111111111),
      .k7(32'b00111101101001010100011100000000),
      .k8(32'b00111101111010010111100010101001),
      .k9(32'b00111100101111101100100100011101)
  ) CON2D_244(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100100010111010100100111),
      .k2(32'b10111101010100111100001101100101),
      .k3(32'b10111101111100111000111100000000),
      .k4(32'b10111100111101100111100111010111),
      .k5(32'b10111110000000011001000110000000),
      .k6(32'b10111100011110110001010111111100),
      .k7(32'b10111011000000111100001001111100),
      .k8(32'b10111011000111010111011011111010),
      .k9(32'b10111101110011100101000110101001)
  ) CON2D_245(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100000100000101111000011010),
      .k2(32'b00111101000101010110000000000111),
      .k3(32'b10111101010000111101001111100011),
      .k4(32'b10111101010110011001010110011111),
      .k5(32'b00111101110011000010000011101100),
      .k6(32'b10111100101011001111011011010000),
      .k7(32'b10111101111010110010101001011000),
      .k8(32'b00111101100100010011111100011001),
      .k9(32'b10111100011011001011001101011101)
  ) CON2D_246(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101101100000001010010010),
      .k2(32'b00111101010100111111110011010101),
      .k3(32'b10111010100110010000111000000011),
      .k4(32'b10111101111100001101010011110111),
      .k5(32'b00111101011010000101100010100001),
      .k6(32'b00111101101100101110100010111110),
      .k7(32'b10111101101000100111100010100000),
      .k8(32'b10111101111010011101011100111011),
      .k9(32'b10111101010011010111011001000110)
  ) CON2D_247(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000110010110001100011100),
      .k2(32'b00111101011111101010101011111010),
      .k3(32'b00111100010101101000010101001001),
      .k4(32'b00111101100111011011011011111110),
      .k5(32'b10111100100111010011001011010010),
      .k6(32'b00111101110110101010110010101010),
      .k7(32'b00111101100101000101010110100011),
      .k8(32'b10111101011100111010101000110001),
      .k9(32'b10111101100100100110111101111110)
  ) CON2D_248(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100001101111011110101101011),
      .k2(32'b00111100100000011010000100011100),
      .k3(32'b10111101110111010110111111101100),
      .k4(32'b00111101000001111100001011111101),
      .k5(32'b00111101000100000010101110101000),
      .k6(32'b10111100110100001010100011011010),
      .k7(32'b00111101010010001011111001001110),
      .k8(32'b10111101000110111110100101010100),
      .k9(32'b00111100110101001010011010010000)
  ) CON2D_249(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010111011000011001100100),
      .k2(32'b10111101111011000000001010011101),
      .k3(32'b00111101110000111111011100101110),
      .k4(32'b10111100111001001110001000010111),
      .k5(32'b00111100100010101110100101010100),
      .k6(32'b00111101100101100111001101110010),
      .k7(32'b00111100010011111111111100011001),
      .k8(32'b00111101001010110100110010111101),
      .k9(32'b10111101010110110011001101110111)
  ) CON2D_250(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001010101001000010101),
      .k2(32'b00111101100100000101001110000111),
      .k3(32'b00111100111010111111010100110001),
      .k4(32'b00111101111001010011111101010011),
      .k5(32'b10111101100111011101111011110000),
      .k6(32'b10111100011010000100111011100000),
      .k7(32'b10111101100010101000011000000111),
      .k8(32'b00111011000101001010001101010101),
      .k9(32'b10111101101100101010001111000101)
  ) CON2D_251(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100010010100001100100101),
      .k2(32'b10111101010110000101000000011111),
      .k3(32'b00111100101011001110001110000010),
      .k4(32'b00111100010011000001100001111010),
      .k5(32'b10111101101001000111110100010000),
      .k6(32'b10111100110111110001111101111100),
      .k7(32'b10111101000110011011010100100111),
      .k8(32'b10111101101111100011001001001110),
      .k9(32'b10111101111110101111011111110100)
  ) CON2D_252(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010101101001111100100010),
      .k2(32'b10111101110111010001100101000001),
      .k3(32'b00111100100010100001100011011001),
      .k4(32'b00111011101100000110100100110101),
      .k5(32'b00111101001011001001011100101100),
      .k6(32'b00111100110110000111010011000111),
      .k7(32'b10111101010110000010011100101001),
      .k8(32'b10111100111110001001001001011010),
      .k9(32'b00111101100011010010110000101101)
  ) CON2D_253(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110010110011110011010011),
      .k2(32'b00111101000101010100110101100110),
      .k3(32'b00111110000000010000111100001000),
      .k4(32'b00111101101000000011101001100100),
      .k5(32'b10111101100111111110010111010101),
      .k6(32'b10111101101111110110110101110000),
      .k7(32'b00111101111101010100110110100111),
      .k8(32'b10111101000010010000010101000010),
      .k9(32'b00111100110101001010000010101011)
  ) CON2D_254(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010101001011100110011010),
      .k2(32'b10111101101100001001110000111100),
      .k3(32'b00111101100011101000010100001011),
      .k4(32'b10111011111011000001011000111110),
      .k5(32'b00111101101110010100000100000100),
      .k6(32'b00111101100000110010110011101000),
      .k7(32'b00111101101110111111110100110111),
      .k8(32'b10111101100010101100001100000001),
      .k9(32'b00111101001001110011001000100011)
  ) CON2D_255(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101010001110001001011000),
      .k2(32'b10111101001110101001111010010011),
      .k3(32'b00111101000100000010111111011011),
      .k4(32'b00111101110100010010000110100101),
      .k5(32'b10111101001001011000110100101001),
      .k6(32'b00111101110000111000100010000011),
      .k7(32'b00111100010000010001000101000010),
      .k8(32'b00111011100000111110000011110101),
      .k9(32'b10111101100001110010001001000100)
  ) CON2D_256(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[15][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011101000110011000000100010)
)   op16(
    .i_pipeline_layer4(i_CORE_IP1[15]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*16-1:DATA_WIDTH*15])
);

/// CON2D_17///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010011001000111001001111),
      .k2(32'b00111101111001010000101011010011),
      .k3(32'b10111101100000011111110110111001),
      .k4(32'b10111101110111001010000010011110),
      .k5(32'b10111101101001010001100011011110),
      .k6(32'b00111100011100111100000011110010),
      .k7(32'b00111101000111011100100110100111),
      .k8(32'b00111101101100110010001011100010),
      .k9(32'b00111101101000101101101011010001)
  ) CON2D_257(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001001100101011000010101),
      .k2(32'b10111101101110101001110101001111),
      .k3(32'b00111011011001000100001000101110),
      .k4(32'b00111101101100011110011011011010),
      .k5(32'b10111101010001000111111000110110),
      .k6(32'b10111101110111100101000000010101),
      .k7(32'b00111101101100001011101110011101),
      .k8(32'b00111100001010111110100001011001),
      .k9(32'b00111101001111100011000000000111)
  ) CON2D_258(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110110000010100100100),
      .k2(32'b00111101001110111100101011110110),
      .k3(32'b00111101101010011000110111100011),
      .k4(32'b00111101100010101101010101111100),
      .k5(32'b00111101010000000100010111100010),
      .k6(32'b00111100010001100100011101101101),
      .k7(32'b00111100100011101100011100101001),
      .k8(32'b00111100100101101111010111001110),
      .k9(32'b00111100110010010111101011110000)
  ) CON2D_259(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101110100011011101100011),
      .k2(32'b00111011110100010011101111001011),
      .k3(32'b00111101000011101100010010110101),
      .k4(32'b10111101010001001010000111001011),
      .k5(32'b10111101001011001111010111101110),
      .k6(32'b10111101100000001011100101011010),
      .k7(32'b10111101101010001011110100111000),
      .k8(32'b00111101101111100000000011010100),
      .k9(32'b00111100110011111111101111000001)
  ) CON2D_260(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100000000000101100101111),
      .k2(32'b10111101101101110111101010001000),
      .k3(32'b10111100001010001011001110101001),
      .k4(32'b10111101111101100101100011011100),
      .k5(32'b10111101101111101011000000011001),
      .k6(32'b00111101011110001111111000100100),
      .k7(32'b00111101110010011010100000110110),
      .k8(32'b10111101110111010111100010001110),
      .k9(32'b10111101110010111111110110100010)
  ) CON2D_261(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011010100010000000010011),
      .k2(32'b00111100111000010001110011010000),
      .k3(32'b10111101101000101101010000011011),
      .k4(32'b00111101010000111110000010111010),
      .k5(32'b00111100100100101110110100101110),
      .k6(32'b00111101101001100000011000101110),
      .k7(32'b00111100010000110001011110101100),
      .k8(32'b10111101101010101011111111110000),
      .k9(32'b00111101101010110100110110001011)
  ) CON2D_262(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011001110101011101100111),
      .k2(32'b00111100110010101101101001101101),
      .k3(32'b10111101100111000111000000011010),
      .k4(32'b00111101001011100011101000000100),
      .k5(32'b00111100001111001100100101010000),
      .k6(32'b10111101001001111110000100100001),
      .k7(32'b10111100111011111110000101001001),
      .k8(32'b00111101101001001010101110000111),
      .k9(32'b10111101101001110001000011101110)
  ) CON2D_263(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100000001011010000110101),
      .k2(32'b00111101111101011011001011100010),
      .k3(32'b00111101011011111101001101001111),
      .k4(32'b00111101010011011011101111110110),
      .k5(32'b00111101010000010011011000101101),
      .k6(32'b00111100111110011010101100001111),
      .k7(32'b00111100111011000000100110011011),
      .k8(32'b10111101110111001010001110001001),
      .k9(32'b10111101011001101000010000100011)
  ) CON2D_264(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101000110101000101111000),
      .k2(32'b00111100111010000101110001111011),
      .k3(32'b10111100101000010001010001111100),
      .k4(32'b10111101100110000100000000101010),
      .k5(32'b10111100110111000000001001110000),
      .k6(32'b00111101100101001101110101010101),
      .k7(32'b00111100011110011011111101000001),
      .k8(32'b10111101000100000101011101101111),
      .k9(32'b10111011100001111001001101101000)
  ) CON2D_265(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010111110111111111011),
      .k2(32'b00111101011010101100101001111101),
      .k3(32'b00111100110100001000111110010101),
      .k4(32'b10111101101000000101110101000111),
      .k5(32'b00111101101111110000111011111011),
      .k6(32'b00111100101100011001101110100001),
      .k7(32'b00111101110100000000001110000000),
      .k8(32'b00111101101001010010110101110010),
      .k9(32'b10111101011111000101001001011011)
  ) CON2D_266(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010000010000011111111011),
      .k2(32'b00111101111100001001111110001000),
      .k3(32'b10111100100010111110010110010100),
      .k4(32'b00111100011001001000000110100101),
      .k5(32'b10111101001110110111010110001010),
      .k6(32'b00111101100101101000110100010001),
      .k7(32'b10111101100000010101100101011110),
      .k8(32'b10111101100110001111110110010010),
      .k9(32'b10111100100011010010100100100111)
  ) CON2D_267(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001001111001111001000101),
      .k2(32'b10111101100101100101101001101100),
      .k3(32'b00111101000101010001000101111010),
      .k4(32'b10111101010000101011111101111100),
      .k5(32'b00111101100000000111111001001011),
      .k6(32'b10111101101011010001100100001000),
      .k7(32'b00111100100111000001001001110010),
      .k8(32'b00111101110000110011000010110111),
      .k9(32'b00111101011100110000001010111001)
  ) CON2D_268(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110101010101010001001111),
      .k2(32'b00111011110110000010110000100010),
      .k3(32'b10111101000010001100001110000001),
      .k4(32'b10111011110000100001010011010100),
      .k5(32'b10111101100011111001110001001110),
      .k6(32'b10111101110010010000000001011100),
      .k7(32'b00111100011010011010010100011110),
      .k8(32'b10111101110011001011011100110010),
      .k9(32'b10111100001001110100110010110011)
  ) CON2D_269(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011100111111111011001100010),
      .k2(32'b00111101101110000111111110000000),
      .k3(32'b10111101101010101011110110101011),
      .k4(32'b00111101011100100000011100111010),
      .k5(32'b00111101111010011001101010010001),
      .k6(32'b10111101000010000010000011110010),
      .k7(32'b00111101001001111000100011000101),
      .k8(32'b10111001111000110011010110110110),
      .k9(32'b10111100000100001001111001011001)
  ) CON2D_270(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010000111100110011100001),
      .k2(32'b10111101011000001101010101101010),
      .k3(32'b10111101001001011001010000000110),
      .k4(32'b00111100011100000001001010111010),
      .k5(32'b10111101100101010000011010011001),
      .k6(32'b00111011111100110011010000100001),
      .k7(32'b00111101101101000100011110110001),
      .k8(32'b00111100110000110110001010011110),
      .k9(32'b00111101111110011110111001101000)
  ) CON2D_271(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011001010000111000000),
      .k2(32'b10111101101000111100011000110101),
      .k3(32'b10111101101111101011000001001010),
      .k4(32'b00111011000101110110010100110010),
      .k5(32'b00111101000000001011101101100101),
      .k6(32'b00111101010001100110100010010000),
      .k7(32'b10111101010110010100101010011011),
      .k8(32'b10111101100111110110000111101010),
      .k9(32'b00111100010011111110011010001101)
  ) CON2D_272(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[16][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011111001111101010000001010)
)   op17(
    .i_pipeline_layer4(i_CORE_IP1[16]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*17-1:DATA_WIDTH*16])
);

/// CON2D_18///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100000011111101100110001),
      .k2(32'b10111101011000010101000111101010),
      .k3(32'b10111101100011110011001100001011),
      .k4(32'b10111100101000101010001110011011),
      .k5(32'b10111101100010100111010111101011),
      .k6(32'b00111101011000000110100001011001),
      .k7(32'b00111011100110111111001001101101),
      .k8(32'b10111101001010111111100111011010),
      .k9(32'b10111101011010011111001011001100)
  ) CON2D_273(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001111100000001100110011),
      .k2(32'b10111101001011100010000101011011),
      .k3(32'b10111101000000101111011111001100),
      .k4(32'b10111101101101110110010011110010),
      .k5(32'b00111101001101110100101100110011),
      .k6(32'b00111101100111011010001111110100),
      .k7(32'b00111101100100010011010010000111),
      .k8(32'b10111011010100011010010110001110),
      .k9(32'b00111101100010100010101111111001)
  ) CON2D_274(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111101010110011111100101),
      .k2(32'b00111101110010111001100111100000),
      .k3(32'b00111100100110100000010110110001),
      .k4(32'b00111101110110100010000111001001),
      .k5(32'b10111101101011010010001001100000),
      .k6(32'b00111101001001101101101101111000),
      .k7(32'b10111101101000100100100100011101),
      .k8(32'b00111101101111011110101010001001),
      .k9(32'b00111101011111101110111101000100)
  ) CON2D_275(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111000000010100101011110),
      .k2(32'b10111101001011000001110010111101),
      .k3(32'b10111000100011111011100101101110),
      .k4(32'b00111101110010100111001100010101),
      .k5(32'b10111101010010001101110011000011),
      .k6(32'b00111101110110010001001000000100),
      .k7(32'b10111101011110101101000101010110),
      .k8(32'b00111101101110101011001101001110),
      .k9(32'b10111011001011001111011000111010)
  ) CON2D_276(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110110011010011110010111),
      .k2(32'b00111101011101011100110100010111),
      .k3(32'b10111100110101001001110111010011),
      .k4(32'b00111011100000010001110001101010),
      .k5(32'b00111101111000000110000000011001),
      .k6(32'b10111101100101000001100000100100),
      .k7(32'b00111101001111110101100100011000),
      .k8(32'b00111101101100011010001011100110),
      .k9(32'b00111101100101110100011010100011)
  ) CON2D_277(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110000101011101000011100),
      .k2(32'b00111101101001100000111110111110),
      .k3(32'b00111100010000001101011000001100),
      .k4(32'b00111100001100000011111001101101),
      .k5(32'b10111100110101111100000000011101),
      .k6(32'b10111101111000001101000110100011),
      .k7(32'b10111101100111010111100110110010),
      .k8(32'b00111101010101100100011011100101),
      .k9(32'b10111101101011001100010001011111)
  ) CON2D_278(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111101101101100010111010),
      .k2(32'b00111101011000000001001000011010),
      .k3(32'b10111101001010011010111101101010),
      .k4(32'b00111101000100011001001101001100),
      .k5(32'b10111101111000111000000001001010),
      .k6(32'b10111100110001111000111100110101),
      .k7(32'b00111101101101111011000001100001),
      .k8(32'b00111101001010111001000000110101),
      .k9(32'b00111101001111111010001001011101)
  ) CON2D_279(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100111000101010010011101),
      .k2(32'b00111101101001001000110011100011),
      .k3(32'b10111100001111111000101000001111),
      .k4(32'b00111101101010100000101010011101),
      .k5(32'b10111100100011111111111101010100),
      .k6(32'b00111101011111110011000100110110),
      .k7(32'b00111101000111100010000000110000),
      .k8(32'b10111101100011010011100111101101),
      .k9(32'b00111101100010111110010001000011)
  ) CON2D_280(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001101001000100011100111),
      .k2(32'b00111101111100000000110010001011),
      .k3(32'b10111101100110100001011011000110),
      .k4(32'b00111101010001011100111010000100),
      .k5(32'b00111101010110011011101001001010),
      .k6(32'b10111101101101100011100000000100),
      .k7(32'b00111101111100010011010100111111),
      .k8(32'b10111101100011111100011000110011),
      .k9(32'b10111101101110001000101011111010)
  ) CON2D_281(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011000011110001101011000),
      .k2(32'b10111101010100000101111100001011),
      .k3(32'b00111101000111101001011001011001),
      .k4(32'b10111101100010111111111100111010),
      .k5(32'b10111101001101011001101101001110),
      .k6(32'b00111101111000010011000000100000),
      .k7(32'b00111100101100000101110110001010),
      .k8(32'b10111101001000110110111000000010),
      .k9(32'b00111101000001000101110101000101)
  ) CON2D_282(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111101110001010001111010),
      .k2(32'b10111100100010111001011111111000),
      .k3(32'b10111101000111010011000001001101),
      .k4(32'b10111101110101010101011110011111),
      .k5(32'b10111101010110101110000010110101),
      .k6(32'b10111101011001110000111111010011),
      .k7(32'b00111101010101000101001100110110),
      .k8(32'b00111100000010010011000100101011),
      .k9(32'b00111101000011011000111010011110)
  ) CON2D_283(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100111101101100110101110),
      .k2(32'b00111101101110101110001101000000),
      .k3(32'b00111101101010110000101101101010),
      .k4(32'b00111101111001110000010001101111),
      .k5(32'b00111101110111101100000011001010),
      .k6(32'b10111101011010100010001011011110),
      .k7(32'b10111101101001011001010101110100),
      .k8(32'b00111101000110111110110101000001),
      .k9(32'b10111101000011001000101001000010)
  ) CON2D_284(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100010110111010111110111),
      .k2(32'b00111101010101010011011000011111),
      .k3(32'b00111101000011001011010111000110),
      .k4(32'b10111101110110000110010100000011),
      .k5(32'b10111101010001001001111110100110),
      .k6(32'b00111101100111001110101101100001),
      .k7(32'b00111101001100111000010110101000),
      .k8(32'b00111010100111100001010111101100),
      .k9(32'b00111101000100011100101010011101)
  ) CON2D_285(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100111101011110010100011),
      .k2(32'b00111011100110111100011011010110),
      .k3(32'b10111101001010100000010011110111),
      .k4(32'b10111100110000010110100000011010),
      .k5(32'b10111101101111010011001111100101),
      .k6(32'b00111101001100001010011001010110),
      .k7(32'b10111101101010001100000011100101),
      .k8(32'b10111101110100110111000100101101),
      .k9(32'b00111101011100110000000111000000)
  ) CON2D_286(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101000001100100101000111),
      .k2(32'b10111101101000010010011111011000),
      .k3(32'b10111101101100010110110010001101),
      .k4(32'b10111101110000110100101111101110),
      .k5(32'b00111100100000000010011001101110),
      .k6(32'b00111101100110010111101100110001),
      .k7(32'b00111101010100010001111001101110),
      .k8(32'b00111101110000111000110101000001),
      .k9(32'b00111101101100100000111010001100)
  ) CON2D_287(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000111111101010111010110),
      .k2(32'b00111101000101110100111110010011),
      .k3(32'b00111101110111101111110001100001),
      .k4(32'b10111101000011111001011010011111),
      .k5(32'b10111101100110011010010011100001),
      .k6(32'b00111101100101010100000110001110),
      .k7(32'b00111101110101000001010001111101),
      .k8(32'b00111101101011111000001000110001),
      .k9(32'b00111101000101011000101100011000)
  ) CON2D_288(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[17][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011011000001111100101110100)
)   op18(
    .i_pipeline_layer4(i_CORE_IP1[17]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*18-1:DATA_WIDTH*17])
);

/// CON2D_19///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010111101111010110111011),
      .k2(32'b00111101110110110001100111101111),
      .k3(32'b00111101101101100000001001001110),
      .k4(32'b10111100010000000011001101011001),
      .k5(32'b10111101101110101111000001101001),
      .k6(32'b00111101111011000110000011101010),
      .k7(32'b10111101111100001000000010100010),
      .k8(32'b00111010100011010010001000101110),
      .k9(32'b00111101100001010100000001110001)
  ) CON2D_289(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010011010011111000001110),
      .k2(32'b10111101101010110111111110000110),
      .k3(32'b00111101111011111000000011000100),
      .k4(32'b00111100011101110110100011011010),
      .k5(32'b10111101100000010000110111011101),
      .k6(32'b10111101100110001010101110010001),
      .k7(32'b00111100111010001110101111101010),
      .k8(32'b00111101111110001001100000001100),
      .k9(32'b00111110000100111100010011101000)
  ) CON2D_290(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111010110100110110100110),
      .k2(32'b00111100010010001100110110000100),
      .k3(32'b00111101111011011110010110111010),
      .k4(32'b00111101100100011000110111110101),
      .k5(32'b00111100001001101001111010010111),
      .k6(32'b10111101101111010101111111101100),
      .k7(32'b00111101000001011010100011010000),
      .k8(32'b00111101110001000010111010111110),
      .k9(32'b10111101111001101110000101111110)
  ) CON2D_291(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010011001101011000010001),
      .k2(32'b00111101011001111100110100001110),
      .k3(32'b00111101110101111011110101000100),
      .k4(32'b10111011110110110101110001010010),
      .k5(32'b00111101101111011100110110001101),
      .k6(32'b00111101000110011101100100111011),
      .k7(32'b10111100100110100111010000110011),
      .k8(32'b00111100100111000010010110110010),
      .k9(32'b00111101110011010110111101100110)
  ) CON2D_292(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110000101111001001110000),
      .k2(32'b00111101011101011100000010011001),
      .k3(32'b00111101111100101000010110101011),
      .k4(32'b00111101000101000110111000000111),
      .k5(32'b00111101110001110101110000101110),
      .k6(32'b00111101001010010100101000101100),
      .k7(32'b00111101000111111001000111111110),
      .k8(32'b00111101101110101010101111000000),
      .k9(32'b00111100100001011011111110101011)
  ) CON2D_293(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100010010101110111111100),
      .k2(32'b00111101000010000010100010011110),
      .k3(32'b10111101101001000111011111100111),
      .k4(32'b00111101111000101100001011001001),
      .k5(32'b10111101110110010010101111011100),
      .k6(32'b00111101011101010100100010100110),
      .k7(32'b00111101100001001011101010111100),
      .k8(32'b10111100101110101011001000101111),
      .k9(32'b10111101101001100000100101011001)
  ) CON2D_294(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100100001100101011010000),
      .k2(32'b10111101100111101111010101110011),
      .k3(32'b00111101001111100010100010010001),
      .k4(32'b00111101010000111010101100001010),
      .k5(32'b00111100011100011010000011001101),
      .k6(32'b00111100001100000111011101001110),
      .k7(32'b00111101110100001000110101010111),
      .k8(32'b10111101101010110010100011100011),
      .k9(32'b10111100111001101010010001111001)
  ) CON2D_295(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100000110010000110110100),
      .k2(32'b10111101000111100000011111000010),
      .k3(32'b00111101110111101000111100111101),
      .k4(32'b10111101000010000110011001100110),
      .k5(32'b10111101010000011000011001100100),
      .k6(32'b00111101100010000001100101100010),
      .k7(32'b00111100011110000111101000110101),
      .k8(32'b10111011111111001110110011001000),
      .k9(32'b10111101110111001101010100100000)
  ) CON2D_296(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101101101011111000001011),
      .k2(32'b10111101100111001000011100101110),
      .k3(32'b00111101011110111100011011010010),
      .k4(32'b00111101110000101110110101000010),
      .k5(32'b10111101010000001001110001111011),
      .k6(32'b00111101000101010100111111010110),
      .k7(32'b00111101011001101111001111000000),
      .k8(32'b10111101100111000011111111001010),
      .k9(32'b00111101100011000100101011110110)
  ) CON2D_297(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011011001000010001011101),
      .k2(32'b10111101110101000100111101100000),
      .k3(32'b10111100011010111110111100001110),
      .k4(32'b10111101101011000011111001100111),
      .k5(32'b00111101100010101111000101110101),
      .k6(32'b00111101111001110011101111100011),
      .k7(32'b10111010110111110010000001010010),
      .k8(32'b00111101101111010010000010011011),
      .k9(32'b10111011011101001101111100000001)
  ) CON2D_298(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001001001111001100010111),
      .k2(32'b00111101110101001010011100010001),
      .k3(32'b10111101100110110010000010100011),
      .k4(32'b10111101111110101101100111000110),
      .k5(32'b10111101100001101110111110010001),
      .k6(32'b00111101010100011101100111011001),
      .k7(32'b00111100101110110101001111000110),
      .k8(32'b10111101101000011000100110010110),
      .k9(32'b10111101101001111010101100111110)
  ) CON2D_299(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100101110110111011110),
      .k2(32'b10111101010110111010100100010000),
      .k3(32'b00111101001011101101000001111000),
      .k4(32'b10111101101110111000101101011101),
      .k5(32'b00111101011001000110101001010110),
      .k6(32'b10111101000100000011100000000001),
      .k7(32'b10111101010011011010110110110001),
      .k8(32'b00111101111000000010100110110000),
      .k9(32'b00111101101000100111000000010010)
  ) CON2D_300(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110011010000101001001111),
      .k2(32'b00111101110111011000000110000001),
      .k3(32'b00111011110001111010111110000111),
      .k4(32'b10111011010010010000101010010110),
      .k5(32'b00111011100101001100100010101100),
      .k6(32'b10111101000100011100010111011101),
      .k7(32'b10111101111000010101101001110011),
      .k8(32'b10111101000010011001001000010011),
      .k9(32'b10111100001000010100101100011010)
  ) CON2D_301(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011011100000110101110010),
      .k2(32'b10111101101110001110011110101000),
      .k3(32'b10111101100011000000111111010110),
      .k4(32'b00111100111111110010000101110110),
      .k5(32'b00111101001111001001110000110010),
      .k6(32'b00111101000000101101010000000010),
      .k7(32'b00111101100101100101110111000101),
      .k8(32'b10111101001100101000111110100001),
      .k9(32'b00111101110110111101110000001111)
  ) CON2D_302(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011000011010011110101101),
      .k2(32'b10111101100111100001110011111101),
      .k3(32'b10111101101000011000011010011110),
      .k4(32'b10111101100011101110110111001111),
      .k5(32'b10111100101011010001110100110100),
      .k6(32'b10111101000111100010100011111110),
      .k7(32'b10111100000100001001000011000101),
      .k8(32'b00111100010001111010000110010111),
      .k9(32'b00111101100000101100111001100001)
  ) CON2D_303(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110000010001111001011011),
      .k2(32'b00111100011100110000111011111110),
      .k3(32'b10111001001001111100111111011101),
      .k4(32'b00111101111111010110101111001110),
      .k5(32'b10111101011001111101011001011110),
      .k6(32'b00111101001101000110011110001101),
      .k7(32'b10111100110011011001100101000100),
      .k8(32'b00111100001001110100011000001001),
      .k9(32'b10111101001111111000101101101110)
  ) CON2D_304(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[18][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011101101111101001111111000)
)   op19(
    .i_pipeline_layer4(i_CORE_IP1[18]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*19-1:DATA_WIDTH*18])
);

/// CON2D_20///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101011110001110010111101),
      .k2(32'b00111010000110100111111010111110),
      .k3(32'b00111101100001111010110010110011),
      .k4(32'b00111101100110101001100110110011),
      .k5(32'b00111101011110001101101100101010),
      .k6(32'b10111100111001001111111111100010),
      .k7(32'b10111101100000000100110111000000),
      .k8(32'b00111100110101110001000010011101),
      .k9(32'b00111100110011010000110000100100)
  ) CON2D_305(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111110000001001110101111),
      .k2(32'b00111101000001011101000101100010),
      .k3(32'b00111100111100110100010111010000),
      .k4(32'b10111100101000101101001110011000),
      .k5(32'b10111101101000001010101010011011),
      .k6(32'b00111101000110110111010001011111),
      .k7(32'b10111101010010000000000110100111),
      .k8(32'b10111011000001100000010110010111),
      .k9(32'b10111101101010000110101010010101)
  ) CON2D_306(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111100000010001010100),
      .k2(32'b10111101110000100100001110010011),
      .k3(32'b00111100111110000001111010111110),
      .k4(32'b10111101100010010111100001100101),
      .k5(32'b00111101010101100010010001000000),
      .k6(32'b00111100011100001000011100111000),
      .k7(32'b10111101100100001101011010111100),
      .k8(32'b10111101010101100011101100000001),
      .k9(32'b00111100100000110110000011001011)
  ) CON2D_307(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110110100010100111011100),
      .k2(32'b00111101010001001100110000000110),
      .k3(32'b00111100100011101101100110100000),
      .k4(32'b00111101000110111011111111010011),
      .k5(32'b10111100110001110111100100001001),
      .k6(32'b00111101001001110100110011110000),
      .k7(32'b00111101100100111101011100111000),
      .k8(32'b10111100100001100110010000011010),
      .k9(32'b10111101100000011010100110110110)
  ) CON2D_308(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011000011010011100010),
      .k2(32'b10111101000110111101000001100011),
      .k3(32'b10111100000110100100000111100010),
      .k4(32'b00111011100100111011010111111010),
      .k5(32'b10111101101011101010111011011100),
      .k6(32'b10111100000110000011011110110110),
      .k7(32'b10111101101110100010100101001110),
      .k8(32'b00111101011111110111100101100101),
      .k9(32'b10111101110110101010111100011010)
  ) CON2D_309(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011110010111101000101010000),
      .k2(32'b10111101000000011110101101110111),
      .k3(32'b10111100010101110011111000101011),
      .k4(32'b10111101101111110111100000011110),
      .k5(32'b00111100100110011100110010111101),
      .k6(32'b10111100100010110101011110010001),
      .k7(32'b00111100111100100110011110111010),
      .k8(32'b10111101101110111001011011111111),
      .k9(32'b00111101101000101000001001110100)
  ) CON2D_310(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000101111111000100101111),
      .k2(32'b10111100101001101010110110111110),
      .k3(32'b00111101101001000110000010000000),
      .k4(32'b10111101000001110101001111000100),
      .k5(32'b00111101010111100101111010001111),
      .k6(32'b00111101000000010000110111101100),
      .k7(32'b10111101110111100110001011010011),
      .k8(32'b00111101100010110001111111110100),
      .k9(32'b10111010101010101100000101001001)
  ) CON2D_311(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101001001000001001011001),
      .k2(32'b00111100110111100100000010100001),
      .k3(32'b00111101010111101010110100110111),
      .k4(32'b10111101110100100001111001010110),
      .k5(32'b00111101100011110101011101000101),
      .k6(32'b00111101111101111111110111110101),
      .k7(32'b10111101110010100100111110001010),
      .k8(32'b00111101100001011101100100011010),
      .k9(32'b10111100110101000111011000111000)
  ) CON2D_312(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111010011101000011111111),
      .k2(32'b00111101100000100000011010011001),
      .k3(32'b00111100100101111010011011101100),
      .k4(32'b00111101110111101000100110000100),
      .k5(32'b10111100111001101010001001000110),
      .k6(32'b10111101101010100010100100000010),
      .k7(32'b00111101011101011101010000000010),
      .k8(32'b10111011111010100101010100001101),
      .k9(32'b10111101101110010000010000110011)
  ) CON2D_313(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111001001100000111110),
      .k2(32'b10111101010101001000000100011101),
      .k3(32'b00111100011111101001001110010111),
      .k4(32'b10111101100010011111000000001001),
      .k5(32'b00111101010101010101011111101000),
      .k6(32'b00111101000100010100010110001111),
      .k7(32'b10111101100111001010110000110101),
      .k8(32'b10111101101100010011100001100111),
      .k9(32'b00111100100001100000100100110111)
  ) CON2D_314(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110011111001111000001100),
      .k2(32'b10111101110101101010110011011010),
      .k3(32'b10111100100101100000000011011011),
      .k4(32'b00111101101001011111010011000100),
      .k5(32'b00111101010000001000111101011100),
      .k6(32'b00111101001010011101011111001011),
      .k7(32'b00111101001110110000100011111000),
      .k8(32'b10111101100110011010000000111111),
      .k9(32'b10111101100010100011111011100001)
  ) CON2D_315(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110100000111110001110101),
      .k2(32'b00111101110100100000000101000110),
      .k3(32'b10111100100011011100110100001011),
      .k4(32'b00111101101000001111111011000100),
      .k5(32'b10111100100100110001001011101011),
      .k6(32'b00111100101101100010111111100110),
      .k7(32'b10111101100010010111100101110100),
      .k8(32'b00111101100101110000010100010001),
      .k9(32'b00111100001101111011010010000100)
  ) CON2D_316(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111111001001000011000),
      .k2(32'b10111100011010101001001101000000),
      .k3(32'b00111101100110101110001000011110),
      .k4(32'b00111101111010001011011101011001),
      .k5(32'b00111101100000011001010100111110),
      .k6(32'b10111100000010111100101001010100),
      .k7(32'b10111100101010111110011000110110),
      .k8(32'b00111101110011001101111100000110),
      .k9(32'b10111101100001111111110111111000)
  ) CON2D_317(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100010011011010001111101101),
      .k2(32'b10111101100101100100001001011000),
      .k3(32'b00111101111001110100011111100111),
      .k4(32'b00111101101010101000011010110000),
      .k5(32'b10111101101010100011111111101110),
      .k6(32'b00111110000000000111010000101001),
      .k7(32'b10111100010010101011111001110111),
      .k8(32'b10111100110111011100110010010001),
      .k9(32'b10111101110011010100111001001101)
  ) CON2D_318(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110011101001011011000),
      .k2(32'b00111101100111101100010001010101),
      .k3(32'b10111101001100100011001101010110),
      .k4(32'b00111101010100101110111101111001),
      .k5(32'b10111101101101100011000011001001),
      .k6(32'b00111101111100000101100001000000),
      .k7(32'b00111101111010000010101011011110),
      .k8(32'b00111101000011010011011000000011),
      .k9(32'b00111011010110110110001001100001)
  ) CON2D_319(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010001111110001111101011),
      .k2(32'b10111101001110001100100001011000),
      .k3(32'b10111101100011001100011011110000),
      .k4(32'b10111101001101000010111010100101),
      .k5(32'b10111101010000001101000101110000),
      .k6(32'b00111100001100011100000010001011),
      .k7(32'b00111010101011100101011010100001),
      .k8(32'b00111101110011000101011001001011),
      .k9(32'b10111101110001110000010000101001)
  ) CON2D_320(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[19][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011110111111000100011110111)
)   op20(
    .i_pipeline_layer4(i_CORE_IP1[19]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*20-1:DATA_WIDTH*19])
);

/// CON2D_21///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110111000011111100001010),
      .k2(32'b10111101100111010001010001010100),
      .k3(32'b10111101110110111110110000001011),
      .k4(32'b10111101101011000101110010110011),
      .k5(32'b00111101011101110111011010111010),
      .k6(32'b10111101100001110000001101010111),
      .k7(32'b10111101100110000111101100111111),
      .k8(32'b10111101011111100010001110000010),
      .k9(32'b10111101100101100011100001110100)
  ) CON2D_321(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010111000011001011110101),
      .k2(32'b00111101101011001011001100000110),
      .k3(32'b00111101111001011000011110110001),
      .k4(32'b10111101101101111101110001001011),
      .k5(32'b00111110000000101100000010101111),
      .k6(32'b00111101000010010110011100000000),
      .k7(32'b00111101100011111010001111001110),
      .k8(32'b00111010101011101000100100110000),
      .k9(32'b10111101100101111111000101001100)
  ) CON2D_322(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111011011001110101110000),
      .k2(32'b10111101000010100100001010010110),
      .k3(32'b10111100110001000010110100101010),
      .k4(32'b00111101101111010000001011100010),
      .k5(32'b00111101100111010110010100100101),
      .k6(32'b00111101101101011111001010000100),
      .k7(32'b00111101101011110101010011000101),
      .k8(32'b00111100110110111010011111000101),
      .k9(32'b00111101010110001100000011010100)
  ) CON2D_323(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101010111011010011100011),
      .k2(32'b00111101100000101001100100000000),
      .k3(32'b10111100110100000100111010010111),
      .k4(32'b00111100001010110100011011011000),
      .k5(32'b00111101000011111111100001001001),
      .k6(32'b00111101110010100001100010010100),
      .k7(32'b10111100100000111010101100001010),
      .k8(32'b00111100111111101000001110000110),
      .k9(32'b00111100101101000100110100001101)
  ) CON2D_324(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101000010110101101010010),
      .k2(32'b00111101100101011101011001011001),
      .k3(32'b10111101110011101101110001011111),
      .k4(32'b00111101100100100011110110101110),
      .k5(32'b10111101111011011101000010000011),
      .k6(32'b10111101110100110110001100100001),
      .k7(32'b10111100100000111110110011110101),
      .k8(32'b10111101101110100100110011000001),
      .k9(32'b00111101010100000001100110100111)
  ) CON2D_325(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011011111100011110000),
      .k2(32'b10111101101101110111100100101111),
      .k3(32'b10111101000001001110001111111001),
      .k4(32'b10111101100101110001100100110010),
      .k5(32'b00111101100110101011110101111100),
      .k6(32'b00111101101101101011101011111010),
      .k7(32'b10111101110100101001010000011000),
      .k8(32'b10111100111001100111011001111011),
      .k9(32'b00111101001011100100001110010100)
  ) CON2D_326(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000010001010101100010111),
      .k2(32'b00111101111101111001111110110011),
      .k3(32'b00111101111001001011010001110100),
      .k4(32'b00111100000001011100100111100011),
      .k5(32'b00111110000100010110001010111101),
      .k6(32'b00111110000000001001000010100010),
      .k7(32'b10111101011111100101001101101000),
      .k8(32'b00111110000000001101110001010111),
      .k9(32'b00111101101001101110101111000001)
  ) CON2D_327(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100101010111100111100011),
      .k2(32'b10111100111111011110001100100101),
      .k3(32'b10111101101001010010110001001101),
      .k4(32'b10111101110000100001011100000011),
      .k5(32'b10111101101011111110100110110011),
      .k6(32'b00111101100101110000001111111010),
      .k7(32'b00111101010010010000010100101111),
      .k8(32'b00111101000001111000100011110000),
      .k9(32'b10111011101101111110011010011000)
  ) CON2D_328(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000001011000101011101000),
      .k2(32'b10111101101111001110001111010000),
      .k3(32'b10111011100001000110001100011001),
      .k4(32'b00111101001011101100100000101011),
      .k5(32'b10111101011111101000110101110000),
      .k6(32'b00111101000011010110000110110010),
      .k7(32'b00111101111001110000101101111011),
      .k8(32'b00111101100011110101100001001110),
      .k9(32'b10111101000000001000110001001011)
  ) CON2D_329(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110111110100010100000111),
      .k2(32'b00111100101100101110000101000110),
      .k3(32'b00111101110100011011001110101100),
      .k4(32'b00111011110101011110101101000101),
      .k5(32'b10111101001100000100000100110011),
      .k6(32'b10111101101100010010111110100110),
      .k7(32'b00111100001011000100000001100100),
      .k8(32'b00111101010110110000101101101101),
      .k9(32'b00111101110010000001011001101111)
  ) CON2D_330(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001011111001010010111),
      .k2(32'b10111101100110101100010010100111),
      .k3(32'b10111101100101000100100100100000),
      .k4(32'b00111110000000110010000100011000),
      .k5(32'b00111101110001011001110111101110),
      .k6(32'b00111100110000110110011011111011),
      .k7(32'b00111101100110010000011000010010),
      .k8(32'b10111011100110110001001011100000),
      .k9(32'b00111101101110111010011001010101)
  ) CON2D_331(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111001011000001011000001000001),
      .k2(32'b10111101010110100011100111011101),
      .k3(32'b00111101100101000001011010100011),
      .k4(32'b00111101110010111010110010111110),
      .k5(32'b10111101100001101110100110110101),
      .k6(32'b10111101001110100011110010011110),
      .k7(32'b10111100111011001010100111100010),
      .k8(32'b00111101111011110111101101011111),
      .k9(32'b10111101011001010100001110110000)
  ) CON2D_332(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110000010001111011110011),
      .k2(32'b10111101010110101011001111100101),
      .k3(32'b00111101111101001100100010110110),
      .k4(32'b10111101010101101110111011100110),
      .k5(32'b00111101111001111110001000101011),
      .k6(32'b00111101101001111110101100101110),
      .k7(32'b10111100100000000010000101010010),
      .k8(32'b10111101000100001000001010111000),
      .k9(32'b10111011111001100001101101011100)
  ) CON2D_333(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000001000100101110101011),
      .k2(32'b10111101010001011100100100110010),
      .k3(32'b00111101000001111111111110110000),
      .k4(32'b10111100000110101011000101110001),
      .k5(32'b10111101101010011000010011010010),
      .k6(32'b10111101011111010110100101000110),
      .k7(32'b10111101001000000011010111110101),
      .k8(32'b10111101000010111010000100011111),
      .k9(32'b10111101100101100111111111111100)
  ) CON2D_334(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110000010100101000001111),
      .k2(32'b00111101101110000001110111111001),
      .k3(32'b00111101110010111110100011100100),
      .k4(32'b10111101011111100111010100011010),
      .k5(32'b10111101010111010110101111110101),
      .k6(32'b00111101100011011110100110010010),
      .k7(32'b00111101111111111100100101011100),
      .k8(32'b10111101001100100111001101001101),
      .k9(32'b00111100101000001111110011101000)
  ) CON2D_335(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111010100100111110000011),
      .k2(32'b00111100110101011100000000110000),
      .k3(32'b10111101010100001010010100001011),
      .k4(32'b00111101100011101100100111101111),
      .k5(32'b00111101000100000100011111001100),
      .k6(32'b00111100110011001100110100110101),
      .k7(32'b10111101011101000101110010001000),
      .k8(32'b10111101100110011111011010001010),
      .k9(32'b00111100101011001100100001100000)
  ) CON2D_336(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[20][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111001101000111100011110010100)
)   op21(
    .i_pipeline_layer4(i_CORE_IP1[20]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*21-1:DATA_WIDTH*20])
);

/// CON2D_22///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100010111011011101101101001),
      .k2(32'b10111101100010011010010001100100),
      .k3(32'b00111101010001000001001110100111),
      .k4(32'b10111100000010001011001010111010),
      .k5(32'b00111101110001100100100110000101),
      .k6(32'b00111101100101001000110101110011),
      .k7(32'b10111100110101001101000110101000),
      .k8(32'b00111101101100011110011001110010),
      .k9(32'b00111101100010000000100011001011)
  ) CON2D_337(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101001110010101111100010),
      .k2(32'b00111101010000001000010101110111),
      .k3(32'b00111101011101110111101001100010),
      .k4(32'b00111101110100111001111101101001),
      .k5(32'b10111101110010001001001110100111),
      .k6(32'b00111011101110101000100100101110),
      .k7(32'b10111101101000010110100000011011),
      .k8(32'b00111101000100010111101000110101),
      .k9(32'b00111100000100110100001101100001)
  ) CON2D_338(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001100111100101110111111),
      .k2(32'b00111100111101010111011000110100),
      .k3(32'b00111101101110110101000010010011),
      .k4(32'b10111101010001100011011101010001),
      .k5(32'b00111101011110010010101011011101),
      .k6(32'b00111100110011110010111000000100),
      .k7(32'b00111101110001111100011111010110),
      .k8(32'b10111101111011100011000001100010),
      .k9(32'b00111101101110101011000101010110)
  ) CON2D_339(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101100011001101101010000),
      .k2(32'b00111101110001101110010111011001),
      .k3(32'b00111110000000111000100000001100),
      .k4(32'b00111100100101110101110000111010),
      .k5(32'b00111101111001111101011001111110),
      .k6(32'b10111101100010110001011111010011),
      .k7(32'b00111101101000110101000000000101),
      .k8(32'b00111100111110010111101010111100),
      .k9(32'b10111101001000100100101101110110)
  ) CON2D_340(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101111011110000010001010),
      .k2(32'b00111101000011011001011101010101),
      .k3(32'b00111101000001111011011101101001),
      .k4(32'b00111100111010010001011100110010),
      .k5(32'b10111100000001110100110100011110),
      .k6(32'b00111100000110101000000000110111),
      .k7(32'b00111101010001110100110101000000),
      .k8(32'b00111100100011000000110000001000),
      .k9(32'b00111101111001101001100101111000)
  ) CON2D_341(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111010100001111111010010000111),
      .k2(32'b00111101100110000010010000100011),
      .k3(32'b10111101101011111001011010101101),
      .k4(32'b00111101001111011011011011001010),
      .k5(32'b10111101110011000111000000000110),
      .k6(32'b00111101001110011111001100001000),
      .k7(32'b10111100101010111110000000110010),
      .k8(32'b10111101101011001100010001111001),
      .k9(32'b00111100010001111111100000001001)
  ) CON2D_342(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100010010011110011110101100),
      .k2(32'b10111100101010110100010100010010),
      .k3(32'b10111101011110101011001011110001),
      .k4(32'b00111100110001100011011110101001),
      .k5(32'b00111100000010100101100110010101),
      .k6(32'b00111101011001101100100001100011),
      .k7(32'b00111101001001011000111111011111),
      .k8(32'b10111101110111100111110101000011),
      .k9(32'b00111101101000110000000111001010)
  ) CON2D_343(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010110111011111100101011),
      .k2(32'b00111101101001110111001010110011),
      .k3(32'b00111101100111101101000010001001),
      .k4(32'b00111101100000101011011100100000),
      .k5(32'b10111100100100011011010011000111),
      .k6(32'b10111011011000100111111100100000),
      .k7(32'b10111101011100110011001111111111),
      .k8(32'b10111101010011111101101000000101),
      .k9(32'b00111101110111001110000100100101)
  ) CON2D_344(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000010100101100110110110),
      .k2(32'b00111101001110011001000110000010),
      .k3(32'b10111101101011011110111011010000),
      .k4(32'b00111101110111010011001100000011),
      .k5(32'b00111101011111100011111101111001),
      .k6(32'b00111101000111001110101010101101),
      .k7(32'b10111101111000001101111001000011),
      .k8(32'b00111100101000101010011110010000),
      .k9(32'b10111100110101111100111110000100)
  ) CON2D_345(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111001110110010100000),
      .k2(32'b00111011101100101001001100000000),
      .k3(32'b00111100001100011111111000010011),
      .k4(32'b00111101111001000101110100010111),
      .k5(32'b00111101011010111010100001100001),
      .k6(32'b00111101110110010001101011000101),
      .k7(32'b00111101101011101111110001011110),
      .k8(32'b00111101110110000001101010101101),
      .k9(32'b00111101101100011010100011111001)
  ) CON2D_346(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101000110010110010110110),
      .k2(32'b10111101111100010010010001110010),
      .k3(32'b00111101111001101110101101101001),
      .k4(32'b10111101101011010110001000000100),
      .k5(32'b00111101110010001011001100011010),
      .k6(32'b10111101100100111010011110011110),
      .k7(32'b00111100010010100101010100000101),
      .k8(32'b00111101100110001101111110000110),
      .k9(32'b10111100101101101011011101011011)
  ) CON2D_347(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011101111100000101100),
      .k2(32'b10111101110101000100010100101110),
      .k3(32'b00111100101001100111011111101011),
      .k4(32'b00111101010011010110011010101010),
      .k5(32'b00111101110010100001000101111000),
      .k6(32'b00111101001001011011011001001000),
      .k7(32'b00111100110101001100100000011111),
      .k8(32'b00111101110101010001011101010011),
      .k9(32'b00111101101110010010011101001110)
  ) CON2D_348(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001000111011110100111101),
      .k2(32'b00111101011111100111011010011100),
      .k3(32'b10111101011011000001010100111101),
      .k4(32'b00111101100110011101111010010000),
      .k5(32'b00111101100001110010011101001101),
      .k6(32'b10111101100111100010000100111100),
      .k7(32'b00111011111111110110001000000001),
      .k8(32'b00111101001000011010011001011100),
      .k9(32'b10111100110000011000001110111011)
  ) CON2D_349(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110000001011011100000001),
      .k2(32'b00111101011010011101011101100100),
      .k3(32'b00111101111100000101101100010101),
      .k4(32'b00111100110101100010001010111110),
      .k5(32'b00111101100110000010000111100011),
      .k6(32'b00111110000011111011010010010101),
      .k7(32'b10111101001100000010000111111100),
      .k8(32'b10111101001001110100010000000110),
      .k9(32'b10111100011000011011110010100000)
  ) CON2D_350(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010110010100111001001101),
      .k2(32'b10111110000001000010001101100111),
      .k3(32'b00111101100110000011101110110110),
      .k4(32'b10111100111010010011101011111111),
      .k5(32'b10111101100111001111101000011001),
      .k6(32'b00111011000101101011000110110000),
      .k7(32'b10111101100111010011111001001110),
      .k8(32'b10111101110101010000100001000100),
      .k9(32'b00111101110100001111010101110111)
  ) CON2D_351(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001110000011011000110010),
      .k2(32'b10111101010101001000011010110001),
      .k3(32'b10111010100010001001010000001101),
      .k4(32'b00111100100110011100110100101111),
      .k5(32'b00111101110001101010111101110000),
      .k6(32'b00111101110011111100110110011001),
      .k7(32'b10111101101001010001100101011100),
      .k8(32'b00111101101100101000111100010110),
      .k9(32'b10111101111000010111100011111010)
  ) CON2D_352(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[21][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011010110010001100001100010)
)   op22(
    .i_pipeline_layer4(i_CORE_IP1[21]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*22-1:DATA_WIDTH*21])
);

/// CON2D_23///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000101111110010011010111),
      .k2(32'b10111101100010101111110111010111),
      .k3(32'b00111101000110100000010011011011),
      .k4(32'b00111100111000111001000010011011),
      .k5(32'b00111101100100000010111010110000),
      .k6(32'b00111011001101101000101111110011),
      .k7(32'b10111101001111011001101000110011),
      .k8(32'b10111101100100011010100010111001),
      .k9(32'b00111101100100011001100101001001)
  ) CON2D_353(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111101111001100101111110),
      .k2(32'b00111101001000111100101001110111),
      .k3(32'b10111101010001011000111001011000),
      .k4(32'b10111101110110011011010001010001),
      .k5(32'b00111101100010011001000001111100),
      .k6(32'b10111101000100011110100111100101),
      .k7(32'b00111101001010110101101100001001),
      .k8(32'b00111101000110001110100101111010),
      .k9(32'b00111100101011011111011101000010)
  ) CON2D_354(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110101001010111010101001),
      .k2(32'b00111101010001100101000111000100),
      .k3(32'b00111100100010001110000101010011),
      .k4(32'b00111101001000010110000100101010),
      .k5(32'b10111101101101110001001110010100),
      .k6(32'b00111101111000101111000001101100),
      .k7(32'b00111101100001110111110101101011),
      .k8(32'b00111101101110010011010101101100),
      .k9(32'b10111101100010110010111011000000)
  ) CON2D_355(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000010001101010101011001),
      .k2(32'b10111101110010001110110100000110),
      .k3(32'b00111101001011110110001001100000),
      .k4(32'b00111011110100001100001010101000),
      .k5(32'b00111101001010011010011110011100),
      .k6(32'b00111011111110100111011011000001),
      .k7(32'b10111101110110011011111001011011),
      .k8(32'b10111101100100010111101010110000),
      .k9(32'b10111101101010000011100001111010)
  ) CON2D_356(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100100101001100000011010),
      .k2(32'b00111101000101110111101111001110),
      .k3(32'b10111101101101010000100010001111),
      .k4(32'b10111101110100010001101100111101),
      .k5(32'b10111101011010000110101101100010),
      .k6(32'b10111101110010010111000100111011),
      .k7(32'b10111101010101101111110000100000),
      .k8(32'b00111101010110001000111010100001),
      .k9(32'b10111101110010100000110101001111)
  ) CON2D_357(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101011000110011101111001),
      .k2(32'b10111100010010100111000000010010),
      .k3(32'b10111101111000101100011110111110),
      .k4(32'b00111101111101100111110001001000),
      .k5(32'b00111101111010010000001000000001),
      .k6(32'b00111100111001101110010110111001),
      .k7(32'b00111101100010010000011110101110),
      .k8(32'b00111101111000001010110101001100),
      .k9(32'b00111011001101111000011010010101)
  ) CON2D_358(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000111111111000011100011),
      .k2(32'b10111101011010111111101101000100),
      .k3(32'b10111101111000011001010001010100),
      .k4(32'b10111101010001011000000010111101),
      .k5(32'b10111101000101000001001010111000),
      .k6(32'b00111101010111100000110011010011),
      .k7(32'b10111101001011001101000010110101),
      .k8(32'b00111101101101111111101101100010),
      .k9(32'b10111101101001011000011100000001)
  ) CON2D_359(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011010000000001000111100),
      .k2(32'b10111101100101100111100111110101),
      .k3(32'b00111101010100100100010100101110),
      .k4(32'b10111101011111110001110011100011),
      .k5(32'b10111101011111010101101110101000),
      .k6(32'b00111101101100110110110110000000),
      .k7(32'b10111101101011110100100000010111),
      .k8(32'b10111101101110101100001110011111),
      .k9(32'b00111011110010101000110010000010)
  ) CON2D_360(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111110101010010110011),
      .k2(32'b00111101100101011011001001111010),
      .k3(32'b00111101101001001011001011111111),
      .k4(32'b10111011101110100001111010001110),
      .k5(32'b00111101111001111101101011111101),
      .k6(32'b00111101000001011001110101001011),
      .k7(32'b10111101000010100011011110001101),
      .k8(32'b10111101001111111011011011101111),
      .k9(32'b00111101100001110011100101101001)
  ) CON2D_361(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111111001101010001000000),
      .k2(32'b10111101101011111010100001110010),
      .k3(32'b00111100101100011100110100001011),
      .k4(32'b00111101111111110110110100101001),
      .k5(32'b10111101110001000001111011110100),
      .k6(32'b10111101100101101000011110010110),
      .k7(32'b00111101011101101111011100010000),
      .k8(32'b00111101011101001001000001101110),
      .k9(32'b10111100110110110001010011111011)
  ) CON2D_362(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111110110111111100100011),
      .k2(32'b10111100011111001100110011100000),
      .k3(32'b00111101110101010111101000110001),
      .k4(32'b00111101010111110001011101111011),
      .k5(32'b10111101100010111011101001011010),
      .k6(32'b00111101110000001001000001110110),
      .k7(32'b10111101100111011101010110101011),
      .k8(32'b10111101110001000111111000011100),
      .k9(32'b00111101000001000110000001100000)
  ) CON2D_363(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100110110000101010011101110),
      .k2(32'b10111101110100001001111101000111),
      .k3(32'b00111101001000011100000111000101),
      .k4(32'b00111101110101101010101100101010),
      .k5(32'b00111101100010110100000100100101),
      .k6(32'b00111101100010000000100011111011),
      .k7(32'b00111101000011110000110011100100),
      .k8(32'b00111101110110111110001001111001),
      .k9(32'b10111101101010000101000001000110)
  ) CON2D_364(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111010001011110111010000),
      .k2(32'b10111101100100100110001110011111),
      .k3(32'b10111101111000010000010010010000),
      .k4(32'b00111101100011010010011000111101),
      .k5(32'b10111100100111101010001101101101),
      .k6(32'b00111101101001101100011111000110),
      .k7(32'b10111101100110001011000111010111),
      .k8(32'b10111101101100100000010101000000),
      .k9(32'b00111101101000000011001001010101)
  ) CON2D_365(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100001110111100000111101),
      .k2(32'b00111101010001011111101000001010),
      .k3(32'b10111011111110000001011100000001),
      .k4(32'b10111100100001100100100111101111),
      .k5(32'b00111011110101101100111111101101),
      .k6(32'b00111100111011010001001011011100),
      .k7(32'b10111100100010011110101001011101),
      .k8(32'b00111011100001011000000110010110),
      .k9(32'b00111011111010111100100010111111)
  ) CON2D_366(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101111110010000001000000),
      .k2(32'b10111101010011101101001111010011),
      .k3(32'b00111101111001011111110111110010),
      .k4(32'b00111100110111110010101100101001),
      .k5(32'b10111101101011111101011111001001),
      .k6(32'b10111100100100000110100001010111),
      .k7(32'b00111101101100100011001110110111),
      .k8(32'b00111101110001010110101010101110),
      .k9(32'b00111101110001111100010010011010)
  ) CON2D_367(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100000100110011000000001110),
      .k2(32'b10111101110010000000110010000101),
      .k3(32'b10111100111001100001110101000011),
      .k4(32'b00111101111001100111011011000000),
      .k5(32'b00111100100101000111100010011100),
      .k6(32'b00111101011010011111001011101010),
      .k7(32'b00111101001111100110011100111101),
      .k8(32'b00111101101010110010010101100010),
      .k9(32'b10111101011111001011000110011110)
  ) CON2D_368(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[22][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100001110000100110101101100)
)   op23(
    .i_pipeline_layer4(i_CORE_IP1[22]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*23-1:DATA_WIDTH*22])
);

/// CON2D_24///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100001101011100110001101010),
      .k2(32'b00111101001000111111100111010101),
      .k3(32'b00111101110000101110111100111001),
      .k4(32'b00111101100001101110001111101110),
      .k5(32'b10111011101010100101101001011100),
      .k6(32'b00111101011101101000101010000011),
      .k7(32'b00111101101010011100001000001011),
      .k8(32'b00111101100111000110111110011000),
      .k9(32'b00111101010110001011000001011000)
  ) CON2D_369(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111010000110010000111100),
      .k2(32'b10111101100011011011010111001100),
      .k3(32'b10111100110010111001001000101111),
      .k4(32'b00111101000011000100101100101000),
      .k5(32'b10111101101111101110001010011001),
      .k6(32'b10111100001001110110101000100011),
      .k7(32'b00111100101001110000110100101011),
      .k8(32'b00111011100010110100101000100001),
      .k9(32'b10111101110110001010001000001111)
  ) CON2D_370(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010001110110101110101001),
      .k2(32'b10111011001101011000001111011100),
      .k3(32'b00111101001100001100001101000100),
      .k4(32'b10111101111011010101111110011100),
      .k5(32'b10111101110110101001000001111001),
      .k6(32'b00111101110010000011011101011110),
      .k7(32'b00111101011110101000011011010111),
      .k8(32'b00111100100111000000001110111000),
      .k9(32'b10111101110011100101010111001100)
  ) CON2D_371(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100110011110011001110011),
      .k2(32'b00111101110010010110100001000000),
      .k3(32'b10111101110111001111000000111101),
      .k4(32'b10111101000000000001101000011111),
      .k5(32'b00111101001010111010001111010001),
      .k6(32'b00111100111010000010011010000111),
      .k7(32'b10111101100000101001011110010100),
      .k8(32'b00111101100011010000010101101100),
      .k9(32'b00111100011000111001001111011110)
  ) CON2D_372(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100011000001011111100111),
      .k2(32'b00111101111100001011100001101111),
      .k3(32'b00111100110000100010110111100110),
      .k4(32'b00111101110101011010100101111101),
      .k5(32'b00111101111000101110010000111111),
      .k6(32'b00111101111010011000001001111111),
      .k7(32'b10111101010000110110011011001001),
      .k8(32'b10111101100011001011001011111110),
      .k9(32'b10111101001111011000110100001011)
  ) CON2D_373(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011000001100010000001010),
      .k2(32'b10111101101110101110101010001000),
      .k3(32'b00111101001001001100001011110000),
      .k4(32'b00111101010000110101000001010111),
      .k5(32'b00111101010000111000100010101100),
      .k6(32'b10111101101001101011011110101001),
      .k7(32'b10111101110000101111010001111010),
      .k8(32'b00111101101001010000001000000111),
      .k9(32'b10111101000100010100101111010001)
  ) CON2D_374(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011101000111010000110110),
      .k2(32'b10111101100100000010011000101101),
      .k3(32'b00111100011101100111001101010110),
      .k4(32'b00111101000100111010010100111110),
      .k5(32'b10111100111010110000110010010110),
      .k6(32'b10111101111011100111110110110000),
      .k7(32'b10111101101001111011101101100111),
      .k8(32'b00111100000100010000010001001100),
      .k9(32'b10111101100101000000110110111001)
  ) CON2D_375(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011100111000000011011),
      .k2(32'b00111100110100110011110101000101),
      .k3(32'b10111100100101110101110011110100),
      .k4(32'b10111101011011010101010000100011),
      .k5(32'b10111100010000010110010100100010),
      .k6(32'b10111101111001011000010000110001),
      .k7(32'b00111101101110000000111100111011),
      .k8(32'b00111101101010100001101001111111),
      .k9(32'b10111101000111001100101011110011)
  ) CON2D_376(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111001100100101010001101),
      .k2(32'b10111011010000110111011111010100),
      .k3(32'b00111101101011100001101000101000),
      .k4(32'b00111101111011100101000101010011),
      .k5(32'b10111011101111011111000101111100),
      .k6(32'b00111101000101010010000101011101),
      .k7(32'b00111100101000010010111000000110),
      .k8(32'b00111100010000101010111001000101),
      .k9(32'b10111100101000111010011010001111)
  ) CON2D_377(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001111011010111111000101),
      .k2(32'b10111101001011000101100111001101),
      .k3(32'b10111101111100001111000101010111),
      .k4(32'b10111101010101111010111001010111),
      .k5(32'b10111101001010001010100000011100),
      .k6(32'b10111101110011001110110111101000),
      .k7(32'b00111101010100011011101011111111),
      .k8(32'b00111101010111000010011000010110),
      .k9(32'b10111100001000110011001011011011)
  ) CON2D_378(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001010011011101100000),
      .k2(32'b10111101111000100111001001101110),
      .k3(32'b10111101011100110100100110010101),
      .k4(32'b00111101000100001001100001101101),
      .k5(32'b00111101101001001100111101011111),
      .k6(32'b00111101101001001110011010011010),
      .k7(32'b00111101101100110001110011101101),
      .k8(32'b10111100011110100101001000010001),
      .k9(32'b00111101110100101110100011010101)
  ) CON2D_379(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110111110011111010101001),
      .k2(32'b10111101100010100000010110101010),
      .k3(32'b10111101100010111000110001010011),
      .k4(32'b00111101001001101110000001000111),
      .k5(32'b10111101011000001011101010010001),
      .k6(32'b00111101101010010101110001101100),
      .k7(32'b10111101011101001111110110010111),
      .k8(32'b10111101100110010010011001010010),
      .k9(32'b00111101101100100001011111011100)
  ) CON2D_380(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011010010001111110110),
      .k2(32'b00111101001101011111110010101000),
      .k3(32'b10111101100111110011111100110011),
      .k4(32'b10111101110110110001110011000011),
      .k5(32'b10111101001001110101101110101010),
      .k6(32'b00111101101101010000000000000001),
      .k7(32'b10111101101111001101110110011001),
      .k8(32'b10111101110111010001000011110110),
      .k9(32'b10111101111100100001111001110110)
  ) CON2D_381(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001100010001110101001),
      .k2(32'b00111101101010010001110101100101),
      .k3(32'b00111101110000000011011101101111),
      .k4(32'b10111101110101000100100000111001),
      .k5(32'b00111101101101000001010111010111),
      .k6(32'b00111101011000001011011101110010),
      .k7(32'b10111101100001101000110010000110),
      .k8(32'b00111100001110111011110110110110),
      .k9(32'b10111011010011110101011101100011)
  ) CON2D_382(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001011101101010000110011),
      .k2(32'b10111100001011000010111101001011),
      .k3(32'b00111100110101111110010110000010),
      .k4(32'b00111101010110000001101110111000),
      .k5(32'b00111101110000001001010000011001),
      .k6(32'b10111110000001011111110000100110),
      .k7(32'b10111011010100010010110001000010),
      .k8(32'b00111101110000110011110000001001),
      .k9(32'b00111101101010001000100011001001)
  ) CON2D_383(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100111100111010100100100),
      .k2(32'b00111101101011010110110010010100),
      .k3(32'b00111101111100000000111101000100),
      .k4(32'b10111101011110101011000111111010),
      .k5(32'b00111101001101100011111010011100),
      .k6(32'b10111011000101001011101001111001),
      .k7(32'b10111101100011111111001001011001),
      .k8(32'b00111101000111001010011011010010),
      .k9(32'b00111100111110100000001011110111)
  ) CON2D_384(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[23][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111010111110000111011000101110)
)   op24(
    .i_pipeline_layer4(i_CORE_IP1[23]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*24-1:DATA_WIDTH*23])
);

/// CON2D_25///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100110110101010111010),
      .k2(32'b00111101101001101010001011011011),
      .k3(32'b00111100010000101111000100101100),
      .k4(32'b00111101101011011110100010100001),
      .k5(32'b00111101110010101101100011011110),
      .k6(32'b10111101101101101010101000001001),
      .k7(32'b10111101111011000001110100000001),
      .k8(32'b10111100100100111100101111110000),
      .k9(32'b10111101110100100011100100000110)
  ) CON2D_385(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010001101110111101110110),
      .k2(32'b10111101110011101111011101111010),
      .k3(32'b00111101101101111101100010000010),
      .k4(32'b10111101100001010011100110000101),
      .k5(32'b00111101100011111111110110111010),
      .k6(32'b10111101001110110011010000001010),
      .k7(32'b10111101010110110011101100010001),
      .k8(32'b00111100001111101001100110000010),
      .k9(32'b10111100101100101011101011000001)
  ) CON2D_386(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001111011111010110111010),
      .k2(32'b00111101100010000010011101011101),
      .k3(32'b00111101111011101010110101001111),
      .k4(32'b00111101110101011011011111111000),
      .k5(32'b00111101111100000011000000000111),
      .k6(32'b10111011111111010101001110010000),
      .k7(32'b00111011110000110111001110110100),
      .k8(32'b00111101110111000101011001101010),
      .k9(32'b00111101011100110010110111100100)
  ) CON2D_387(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100010101001100001001110110),
      .k2(32'b10111101010010001101101010010111),
      .k3(32'b00111101100011100010000101011001),
      .k4(32'b10111010101000111101101110101001),
      .k5(32'b00111101101111000100010000010010),
      .k6(32'b00111101100101011000110011111011),
      .k7(32'b00111100001111011000100000101001),
      .k8(32'b00111101100001101011110100101001),
      .k9(32'b10111101110111010011100000100100)
  ) CON2D_388(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010011100011111011011100),
      .k2(32'b00111101000110110101011111101100),
      .k3(32'b00111101010011101101011101010011),
      .k4(32'b10111100000011000110100001111000),
      .k5(32'b10111101110100111010101001111101),
      .k6(32'b10111011101010110010011110111001),
      .k7(32'b10111101110000100110110010111001),
      .k8(32'b10111101110100010010110011100101),
      .k9(32'b10111101001100001100100100010010)
  ) CON2D_389(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100111011001010100011100),
      .k2(32'b00111101110010000001100011101100),
      .k3(32'b00111101110101110000100100000010),
      .k4(32'b10111011111010101100101100100110),
      .k5(32'b10111101010100111100100010101110),
      .k6(32'b10111100100010110000100010100100),
      .k7(32'b10111101110010000110110100001111),
      .k8(32'b00111101010010001100101111101111),
      .k9(32'b10111101011110001010111001001000)
  ) CON2D_390(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011010010110001110101100),
      .k2(32'b10111101110101111010101111010011),
      .k3(32'b10111101111100000000010111010100),
      .k4(32'b00111101100000001001000110000110),
      .k5(32'b10111101100001111001110100111111),
      .k6(32'b10111101001000000101000110001010),
      .k7(32'b00111100100111110100000110001111),
      .k8(32'b10111101111110111010100111000011),
      .k9(32'b10111010110100100001010000010011)
  ) CON2D_391(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111010101011010010011001),
      .k2(32'b00111101100111110001000011110001),
      .k3(32'b10111000101111101010111110101110),
      .k4(32'b10111011101111001010100100110010),
      .k5(32'b10111101100000001011000001100101),
      .k6(32'b10111101000101110101100101000010),
      .k7(32'b00111101011101001110111010100100),
      .k8(32'b10111101100111110011010100000111),
      .k9(32'b10111100000101011100011011111101)
  ) CON2D_392(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101101000111001011001001),
      .k2(32'b10111101100011100100110100110010),
      .k3(32'b10111101000010011111010001101001),
      .k4(32'b10111101110100000101000001010011),
      .k5(32'b10111101100001110010101110001010),
      .k6(32'b00111101100111100101100010000010),
      .k7(32'b00111101000010010110110111100000),
      .k8(32'b00111101110011111101001011000100),
      .k9(32'b10111100011011001101010001110001)
  ) CON2D_393(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101111011110010000111000),
      .k2(32'b10111101001111000010110000111100),
      .k3(32'b00111101010000010100101011101100),
      .k4(32'b10111101110111011001100110110101),
      .k5(32'b10111100101010101011101101011001),
      .k6(32'b10111100101110010011110011111010),
      .k7(32'b10111101011010111000010011110100),
      .k8(32'b10111101001100000100001101000101),
      .k9(32'b10111101100010110100001111000101)
  ) CON2D_394(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010000000110000001110011),
      .k2(32'b10111100100010110000011100000000),
      .k3(32'b00111101000111011111110001001001),
      .k4(32'b10111101110100001110000010010101),
      .k5(32'b10111100110101001011110101100100),
      .k6(32'b00111101111110001101101011011100),
      .k7(32'b00111101001001000110010110000111),
      .k8(32'b10111101101111110001111110011000),
      .k9(32'b00111100110110001100001101001001)
  ) CON2D_395(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100001110100110111001111),
      .k2(32'b00111101101011100110011000001100),
      .k3(32'b10111101101110010000101101010010),
      .k4(32'b10111100110001001111000101011110),
      .k5(32'b10111101100010100000100011101101),
      .k6(32'b00111101110111001101011010110001),
      .k7(32'b00111011010100001101100110011011),
      .k8(32'b00111100110101100100000100101000),
      .k9(32'b00111101110011100110101111101100)
  ) CON2D_396(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100101001001101000000100),
      .k2(32'b00111100010001100010000110011000),
      .k3(32'b10111101101011000111010101111110),
      .k4(32'b00111101011011000010110001110011),
      .k5(32'b10111011011000001101011111101111),
      .k6(32'b00111101011010011010101000110010),
      .k7(32'b00111101010111100011010010000011),
      .k8(32'b10111100101110110000100110011011),
      .k9(32'b10111101101001011111111010110010)
  ) CON2D_397(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100001010111011010100101),
      .k2(32'b10111100011001011000011100101110),
      .k3(32'b00111101000000100001100101000001),
      .k4(32'b00111101111111010001110011100101),
      .k5(32'b10111101101000100001100010111100),
      .k6(32'b00111101111101000110101011011101),
      .k7(32'b10111011101000100110100010010100),
      .k8(32'b10111011101001111110100011011111),
      .k9(32'b00111100010111100010000000011010)
  ) CON2D_398(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011011111101111001101011),
      .k2(32'b10111100011011001010111110011000),
      .k3(32'b00111101100110011001110110011011),
      .k4(32'b10111011011111001000011010110101),
      .k5(32'b00111101011010010100010110100001),
      .k6(32'b10111101100011111011100001101000),
      .k7(32'b10111101101011011001000110110001),
      .k8(32'b00111101000001100010011000010001),
      .k9(32'b10111101110010110001010001100111)
  ) CON2D_399(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100001011011111000001001),
      .k2(32'b00111101111011001011100111010101),
      .k3(32'b10111101111001011110100111001000),
      .k4(32'b10111101110100010011000000011000),
      .k5(32'b00111100110011100011001110001101),
      .k6(32'b10111101110111111100111110000000),
      .k7(32'b00111101111111110100111110011010),
      .k8(32'b10111101011000110101111011111001),
      .k9(32'b00111101111000111111111011011011)
  ) CON2D_400(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[24][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011100001100000011010001100)
)   op25(
    .i_pipeline_layer4(i_CORE_IP1[24]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*25-1:DATA_WIDTH*24])
);

/// CON2D_26///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110101100101100000111010),
      .k2(32'b10111100111000011110010111011111),
      .k3(32'b00111101111100111011110010010111),
      .k4(32'b00111100101010100000111111011100),
      .k5(32'b00111101001010000010000011011001),
      .k6(32'b10111100110111011101000100010110),
      .k7(32'b00111101110100011111101001001100),
      .k8(32'b00111101110000001101011101101110),
      .k9(32'b00111101100011000001101011001110)
  ) CON2D_401(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111000110000110011001001),
      .k2(32'b10111101101001001100101010110101),
      .k3(32'b10111101000000111001111001101110),
      .k4(32'b10111100110011011111111110011110),
      .k5(32'b10111101101100111011101000100110),
      .k6(32'b00111101111110000001100001000101),
      .k7(32'b00111101000000101001111111001010),
      .k8(32'b00111100101111101010100011010000),
      .k9(32'b10111101011001110100110011011010)
  ) CON2D_402(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011111010010101011001111),
      .k2(32'b00111100101001101001111101101111),
      .k3(32'b00111100000110101101101011111000),
      .k4(32'b10111101110110010010001101000101),
      .k5(32'b10111101100001111100000110000000),
      .k6(32'b10111101110110111010100111100000),
      .k7(32'b10111101100011011010011011111010),
      .k8(32'b10111101100010101101000001111001),
      .k9(32'b00111100110000011001101111100001)
  ) CON2D_403(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011100011100011110101),
      .k2(32'b00111100110110010111001110100001),
      .k3(32'b00111101100000001101011101111011),
      .k4(32'b00111011100110011000100100110010),
      .k5(32'b10111101011010110001000101010010),
      .k6(32'b00111101100100101101110110110011),
      .k7(32'b10111011111001100000000000111110),
      .k8(32'b00111011111011111000100010111010),
      .k9(32'b10111101001110110110100010001101)
  ) CON2D_404(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100110000101010111111100),
      .k2(32'b10111101001001100101101011101000),
      .k3(32'b00111100001000100110100101011000),
      .k4(32'b10111101010111110111010101010101),
      .k5(32'b10111010011100100101111010001100),
      .k6(32'b00111101101001111101001001010100),
      .k7(32'b00111110000000001001001101011101),
      .k8(32'b00111100011100000111100111011110),
      .k9(32'b10111100011111111000110100011011)
  ) CON2D_405(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111001101111100000010010),
      .k2(32'b00111101001111000110010001011001),
      .k3(32'b10111101101110010110011000111001),
      .k4(32'b10111101010110011111100000111000),
      .k5(32'b00111101110000001000010001011111),
      .k6(32'b00111101111000010101000001000011),
      .k7(32'b00111101100111000010000000101011),
      .k8(32'b10111101001100100010111011000100),
      .k9(32'b10111101111011011100110101110001)
  ) CON2D_406(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100101011010010111000100110),
      .k2(32'b00111101001100001101100010111111),
      .k3(32'b00111100110110100000001000011110),
      .k4(32'b10111100111100100100111111000100),
      .k5(32'b00111101100100101110100100011111),
      .k6(32'b10111101001001000101110110101100),
      .k7(32'b10111101101101001101011001100110),
      .k8(32'b00111100010011101000001101111010),
      .k9(32'b10111011001001111110001101100110)
  ) CON2D_407(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011101111101100111001),
      .k2(32'b10111100101111111010101110011100),
      .k3(32'b10111101101100000100101011110111),
      .k4(32'b00111101101001101100100100101100),
      .k5(32'b00111101100101010000111000111000),
      .k6(32'b10111100011100100011010001011010),
      .k7(32'b00111010100000000110010010111000),
      .k8(32'b00111101000000111110100110100110),
      .k9(32'b00111101100100110001001000100110)
  ) CON2D_408(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111010100100000001001010),
      .k2(32'b10111010110110001111001100011101),
      .k3(32'b10111101010100001010010101011010),
      .k4(32'b00111101011010001111001101001001),
      .k5(32'b10111101111100101100001001111100),
      .k6(32'b10111101110100000011101111100110),
      .k7(32'b00111101100111101100010100001110),
      .k8(32'b10111101000010111111000101100110),
      .k9(32'b10111101111011011001100100010110)
  ) CON2D_409(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111110000110110000010001),
      .k2(32'b10111101110011111000011101101011),
      .k3(32'b10111101110010110100110000000100),
      .k4(32'b00111101101111010000001111010000),
      .k5(32'b00111101010100001110001101111111),
      .k6(32'b10111101110110010111011110110101),
      .k7(32'b10111101000111010001000100001111),
      .k8(32'b00111101101010110011101101111110),
      .k9(32'b10111100000010000000100011010110)
  ) CON2D_410(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110011011110000010100110),
      .k2(32'b10111101110101111010100011000010),
      .k3(32'b00111101101001100101010011001110),
      .k4(32'b10111101101111101010000010000011),
      .k5(32'b10111101100000111000100111010000),
      .k6(32'b10111101101100010100000111011101),
      .k7(32'b00111101000110111110100010111101),
      .k8(32'b10111100010000000000110011001110),
      .k9(32'b10111101000001101110100011100011)
  ) CON2D_411(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110101000100111001011111),
      .k2(32'b00111101111111101000101110101011),
      .k3(32'b10111101110100110000001111001001),
      .k4(32'b00111100100101010101111010010001),
      .k5(32'b00111101111010111010110011110000),
      .k6(32'b00111101101101101010010110111101),
      .k7(32'b10111100100100001010111001001011),
      .k8(32'b10111101100011111011100000100000),
      .k9(32'b00111100101010110010010010110111)
  ) CON2D_412(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101100000110001101111000),
      .k2(32'b10111101010101011011100111001101),
      .k3(32'b00111101100010011100011011001110),
      .k4(32'b00111101010011101001111000011000),
      .k5(32'b10111101111001011011001110011010),
      .k6(32'b10111100101110000001111010110110),
      .k7(32'b00111101110010010011010101011111),
      .k8(32'b10111101110110001000110100001111),
      .k9(32'b00111101100100010100011011011111)
  ) CON2D_413(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101011111111011001110011),
      .k2(32'b10111011100100011001010100101101),
      .k3(32'b00111101110000001101001011000000),
      .k4(32'b00111101101001010110111111111000),
      .k5(32'b10111011110111010000100000001101),
      .k6(32'b00111011110100110100100001010001),
      .k7(32'b10111101001101101110010100110010),
      .k8(32'b00111110000011010110101111001000),
      .k9(32'b00111100111100111001101110010010)
  ) CON2D_414(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011101110100010001001100),
      .k2(32'b10111110000000011010100100101111),
      .k3(32'b10111101110011010001011110010110),
      .k4(32'b10111110000001000101011010011110),
      .k5(32'b10111101100010010011001001100101),
      .k6(32'b00111100110010000010111001111111),
      .k7(32'b00111101101101000110000101011110),
      .k8(32'b00111101100100100101111100100001),
      .k9(32'b00111101101110000010001001101110)
  ) CON2D_415(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110100101101111010001),
      .k2(32'b00111101110000100110101100011110),
      .k3(32'b10111101001000010100011100110110),
      .k4(32'b00111101001000011001001011100110),
      .k5(32'b00111101100110101001101011111001),
      .k6(32'b10111100010001010100010101110100),
      .k7(32'b00111101001110111100100010010001),
      .k8(32'b10111101101101110000101111000000),
      .k9(32'b00111011110010011001010011111100)
  ) CON2D_416(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[25][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111011101101010010110111010110)
)   op26(
    .i_pipeline_layer4(i_CORE_IP1[25]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*26-1:DATA_WIDTH*25])
);

/// CON2D_27///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100101000101001101001110100),
      .k2(32'b00111101101001010100110111110111),
      .k3(32'b10111100111110000011000001111000),
      .k4(32'b00111101111100000110010010111110),
      .k5(32'b00111101100111111001111111111111),
      .k6(32'b10111101111000111111100101111001),
      .k7(32'b10111101000111101010010010111111),
      .k8(32'b00111101110101110110110001101010),
      .k9(32'b00111100000101111010000100000110)
  ) CON2D_417(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100010010000010011111110),
      .k2(32'b10111101110110111100100010001001),
      .k3(32'b10111101111000110100001100011111),
      .k4(32'b00111011010011001011100011011011),
      .k5(32'b00111101100010010110111110001000),
      .k6(32'b10111011001010010000011110100011),
      .k7(32'b00111100111100011001110010000000),
      .k8(32'b00111101101110111111000110011101),
      .k9(32'b00111101100000011000000010001110)
  ) CON2D_418(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100111001101001011011011),
      .k2(32'b10111100111010010000100000001111),
      .k3(32'b00111100100001001111011110001111),
      .k4(32'b00111100100101001011000100110000),
      .k5(32'b10111101101100101011110011101001),
      .k6(32'b10111101010000010100110111000101),
      .k7(32'b00111101110000111101001011110111),
      .k8(32'b10111101110101001111111001001000),
      .k9(32'b00111011101110111101111111010100)
  ) CON2D_419(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100010000111000010110010),
      .k2(32'b00111101110100110101011000110011),
      .k3(32'b10111101100100110000101001000100),
      .k4(32'b00111101011110111110100111010011),
      .k5(32'b00111101101010001110110011000010),
      .k6(32'b10111100100110001110100100001010),
      .k7(32'b00111101111101001110111111011011),
      .k8(32'b00111101111101001001100110001110),
      .k9(32'b00111101100111101110010110110011)
  ) CON2D_420(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011011000101011100110000),
      .k2(32'b10111101011011010100100100100000),
      .k3(32'b10111011111011110011000010111110),
      .k4(32'b10111101101001010111111101010010),
      .k5(32'b00111100101101110101111010011011),
      .k6(32'b10111101111000010110001000101000),
      .k7(32'b10111100011110001101001001101011),
      .k8(32'b10111101001000101100010001110011),
      .k9(32'b00111011100111101111011011011110)
  ) CON2D_421(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101101011110011111000101),
      .k2(32'b00111101100001100101100000001011),
      .k3(32'b00111101110000010100000101000000),
      .k4(32'b00111101110100101010011110011001),
      .k5(32'b00111101100000000101011010011011),
      .k6(32'b10111101011110110010111101010110),
      .k7(32'b00111100011100001110011100110100),
      .k8(32'b00111010111010111000001011110010),
      .k9(32'b10111101110110100011010010010001)
  ) CON2D_422(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001001100000010000010100),
      .k2(32'b00111100001110100000111111011100),
      .k3(32'b10111100010110110100101100101110),
      .k4(32'b10111101111110101000011110100110),
      .k5(32'b10111011010011111100100110010111),
      .k6(32'b10111101101011111010000011101011),
      .k7(32'b00111100100010111100001010111101),
      .k8(32'b00111100010111001001000101001010),
      .k9(32'b10111101100011101000001110001000)
  ) CON2D_423(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100000001001001110000011),
      .k2(32'b10111101011011100011000010111101),
      .k3(32'b00111101111010100100101111001101),
      .k4(32'b00111011110001000110010011011010),
      .k5(32'b00111101010100001001001100000110),
      .k6(32'b10111100000100010111100101101000),
      .k7(32'b10111011110101010111111011110111),
      .k8(32'b10111101101110110111110001010110),
      .k9(32'b10111101101000100010101101010010)
  ) CON2D_424(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100000111000111001010),
      .k2(32'b10111101010110011101011110000010),
      .k3(32'b00111101110010000010100001110000),
      .k4(32'b10111100100000101111001000101010),
      .k5(32'b10111101101010101110000001010101),
      .k6(32'b00111101110001010111110111010110),
      .k7(32'b10111101110010101111000100010110),
      .k8(32'b10111101111011111001110000100000),
      .k9(32'b00111101100100010011000110011001)
  ) CON2D_425(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111101010101001001011111),
      .k2(32'b10111101101101000000011000111011),
      .k3(32'b00111101000101101111011000000100),
      .k4(32'b00111100011001100111011011010001),
      .k5(32'b00111101000110110000111001001100),
      .k6(32'b00111101111100011101010111100101),
      .k7(32'b00111101100000111000000010110001),
      .k8(32'b10111101110011110010011001101010),
      .k9(32'b00111101100010010101110100101000)
  ) CON2D_426(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100110101110101101111001),
      .k2(32'b10111101111000001100000110011001),
      .k3(32'b00111101110011010011100111000100),
      .k4(32'b00111100100011000111001110010111),
      .k5(32'b00111101101001011000001101001100),
      .k6(32'b00111101101000101101100100010100),
      .k7(32'b10111101101111001101000000010000),
      .k8(32'b10111101101001001011111110110110),
      .k9(32'b00111101000011001000111110000110)
  ) CON2D_427(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111010101100000101100011001110),
      .k2(32'b00111101010100111010000011111011),
      .k3(32'b10111100000100011101110100110001),
      .k4(32'b10111101001010011110011010000101),
      .k5(32'b10111101001100101010101010011001),
      .k6(32'b00111101110001110000111010111010),
      .k7(32'b10111100101011000101010011101010),
      .k8(32'b10111101100010001101101110000100),
      .k9(32'b00111101110000011110111111000000)
  ) CON2D_428(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101011001101101111011000),
      .k2(32'b10111101100010110010110000011101),
      .k3(32'b00111100111011011011001101000000),
      .k4(32'b00111101100111001000010101001010),
      .k5(32'b10111101011110010011110100010011),
      .k6(32'b00111101010000010011001100100010),
      .k7(32'b10111101011010100110101010000110),
      .k8(32'b10111101010110001101001110111111),
      .k9(32'b10111100010100100101010000101111)
  ) CON2D_429(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111110101101111011101011),
      .k2(32'b00111101001100000100111100110110),
      .k3(32'b10111101011000000100110110010010),
      .k4(32'b10111100011001101111101100110010),
      .k5(32'b00111101011111001010100110000011),
      .k6(32'b10111100001100110111010010101111),
      .k7(32'b00111101101001101010100000110011),
      .k8(32'b00111101111110011001010110100011),
      .k9(32'b00111101010101001001100011011110)
  ) CON2D_430(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100000110100101011000011),
      .k2(32'b00111101011101001011111101000000),
      .k3(32'b00111101101101111011011001000010),
      .k4(32'b10111101101011010111001101010110),
      .k5(32'b00111110000000101010110011111010),
      .k6(32'b00111100100100111111000111011000),
      .k7(32'b00111101000011100101001111000010),
      .k8(32'b00111101000100100100100011111010),
      .k9(32'b10111101011001011100101100011001)
  ) CON2D_431(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100111011001000111010010),
      .k2(32'b10111101000100111101000011111000),
      .k3(32'b00111101100000111011010110000001),
      .k4(32'b00111101110101101100001000111101),
      .k5(32'b00111011100100011010100010110111),
      .k6(32'b10111101101011011010011010111010),
      .k7(32'b10111101011101100100010011001000),
      .k8(32'b10111101100011110001101100101011),
      .k9(32'b10111100111001100000101010010111)
  ) CON2D_432(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[26][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111011100110110101000110100100)
)   op27(
    .i_pipeline_layer4(i_CORE_IP1[26]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*27-1:DATA_WIDTH*26])
);

/// CON2D_28///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111010101011001000111010),
      .k2(32'b10111101011110111100011111110000),
      .k3(32'b00111100100100010001000011001111),
      .k4(32'b10111100100100000110011000010011),
      .k5(32'b10111101101001010100010110110110),
      .k6(32'b00111100101100011001110100100001),
      .k7(32'b00111101010100100110101101001000),
      .k8(32'b00111101010011111111110000100010),
      .k9(32'b10111101111011100000100000011000)
  ) CON2D_433(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101110000000001010000111),
      .k2(32'b10111101000100111101010010101101),
      .k3(32'b10111100111110110101000101101111),
      .k4(32'b10111110000000001011100110110110),
      .k5(32'b00111100100010101110000011100000),
      .k6(32'b10111101011001000010100001000100),
      .k7(32'b00111101101110011001101101110010),
      .k8(32'b10111101001100111000100001001000),
      .k9(32'b00111101110110011001000111111110)
  ) CON2D_434(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111110000000000101101100111111),
      .k2(32'b00111101011101101111111001101110),
      .k3(32'b10111101111111011100011110101000),
      .k4(32'b10111101000100001100110110010110),
      .k5(32'b10111101011100001101010011100001),
      .k6(32'b00111100100010011111111101101001),
      .k7(32'b00111100111001101011111011000011),
      .k8(32'b10111101010111001101011000101111),
      .k9(32'b00111101101101010100011000110001)
  ) CON2D_435(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011001111101111011101100),
      .k2(32'b00111101111000010011101110000001),
      .k3(32'b00111101011000110010100111100010),
      .k4(32'b10111100111110011101100101100111),
      .k5(32'b10111100110110011100001001111110),
      .k6(32'b10111101101101011011001101111011),
      .k7(32'b10111100110011101110110010100011),
      .k8(32'b10111101100100010000101111100011),
      .k9(32'b10111101110100111001100001100111)
  ) CON2D_436(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011100010000111100110111),
      .k2(32'b10111101100010001011100001010101),
      .k3(32'b00111100111011111110011111101110),
      .k4(32'b10111101001100000111100100001111),
      .k5(32'b10111100100000100011100100001110),
      .k6(32'b10111011100101100000101100100001),
      .k7(32'b00111101000011011000001000000010),
      .k8(32'b00111101011001101101101011100100),
      .k9(32'b00111011110000010110111111100010)
  ) CON2D_437(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001110000011000110001000),
      .k2(32'b10111100100000100010111000101011),
      .k3(32'b00111101110001000100111100001001),
      .k4(32'b00111011110100000100100101101010),
      .k5(32'b10111101010111000110010011011111),
      .k6(32'b10111101100110100000110100010011),
      .k7(32'b00111101001000111001101010010111),
      .k8(32'b10111010110011111001110010110101),
      .k9(32'b00111100100101000000010110001010)
  ) CON2D_438(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101010000000100000011100101),
      .k2(32'b00111101100110111011111100000011),
      .k3(32'b00111100000011000011110100110101),
      .k4(32'b00111100110110011001101100010000),
      .k5(32'b10111101101001000000110101110111),
      .k6(32'b10111100101011100110111110000000),
      .k7(32'b10111100110001100110000000000101),
      .k8(32'b10111100011100011011010101001011),
      .k9(32'b00111101011011100101001100010110)
  ) CON2D_439(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011010000000110010110100),
      .k2(32'b00111101110101100100001011111010),
      .k3(32'b10111101011101100011000100010010),
      .k4(32'b00111101110001111000110000100001),
      .k5(32'b00111101110100100010101000100011),
      .k6(32'b00111101101010000101010111101010),
      .k7(32'b00111101100110110100111111101111),
      .k8(32'b00111101100001101000101110101100),
      .k9(32'b10111100100101010110000010010101)
  ) CON2D_440(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100100101010011000011000),
      .k2(32'b10111100110010110110001000110001),
      .k3(32'b10111101110011111011001001000001),
      .k4(32'b10111100001011110110100110011111),
      .k5(32'b00111101000000101101111110111010),
      .k6(32'b00111101101011110001011000111110),
      .k7(32'b10111110000000000011011000111011),
      .k8(32'b10111011111110110000110101001001),
      .k9(32'b10111101100100101111111100111111)
  ) CON2D_441(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011110101010100011000111),
      .k2(32'b00111101000100110111010100010101),
      .k3(32'b10111100101101010111100000010010),
      .k4(32'b10111101001011101100101101011010),
      .k5(32'b00111100111001010100011111010000),
      .k6(32'b10111101101000111101111101011000),
      .k7(32'b00111101101010100110010110100010),
      .k8(32'b10111100110111111110010100000001),
      .k9(32'b10111101100001000101001001110010)
  ) CON2D_442(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010111101100001000000),
      .k2(32'b00111101111010100101110101011110),
      .k3(32'b10111101000101011110001101010100),
      .k4(32'b10111100101101111101001100111110),
      .k5(32'b10111011100110000000111000000011),
      .k6(32'b00111101111100101111100100010110),
      .k7(32'b10111101000010011111011001010101),
      .k8(32'b10111101011010011110101000010100),
      .k9(32'b00111101100111011011010111000101)
  ) CON2D_443(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100011000110100000110100),
      .k2(32'b10111101010111101110100110100000),
      .k3(32'b00111101110000000010100010110110),
      .k4(32'b00111101011101100011001001110010),
      .k5(32'b10111100110101001011110101100101),
      .k6(32'b10111101101000110111101001110110),
      .k7(32'b10111100110001110100001101111000),
      .k8(32'b10111101011100010001111000111111),
      .k9(32'b10111100101000101100100000111111)
  ) CON2D_444(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011001110010101101110100010),
      .k2(32'b00111011111011001101101100011000),
      .k3(32'b00111100100011011011111100000101),
      .k4(32'b10111101110011110101101101100000),
      .k5(32'b00111101101000011110110110100110),
      .k6(32'b10111101000111001001101110111001),
      .k7(32'b10111100000001011111100001000000),
      .k8(32'b10111101010000000001110000100100),
      .k9(32'b00111100110010110001110111001101)
  ) CON2D_445(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001100101000101110000100),
      .k2(32'b00111100111010100100011111101101),
      .k3(32'b00111011110101000011100011110001),
      .k4(32'b00111101100101000111101110111111),
      .k5(32'b10111010001101111001101011001100),
      .k6(32'b00111101000100000100100011011101),
      .k7(32'b00111100110011110010110100010011),
      .k8(32'b10111100110110100011011111001101),
      .k9(32'b10111101011100000011011000011111)
  ) CON2D_446(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110100000110111000001001),
      .k2(32'b00111100000100011110110101000110),
      .k3(32'b00111101010100110000000111001100),
      .k4(32'b10111101001000001001001111010110),
      .k5(32'b00111101011101111100111111101110),
      .k6(32'b10111101100100111001001100101010),
      .k7(32'b00111100101000101110100001011010),
      .k8(32'b10111101100000101001011010111111),
      .k9(32'b10111101101011101101011110101111)
  ) CON2D_447(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011100010111111110110100),
      .k2(32'b10111100010011101101111000011101),
      .k3(32'b00111101100000101100011100111100),
      .k4(32'b10111101110000011101110010100111),
      .k5(32'b10111101001011101100011110111110),
      .k6(32'b00111101001010011110101001010110),
      .k7(32'b10111101100101100010110011101000),
      .k8(32'b10111101111000100110111111001101),
      .k9(32'b10111100100001110101101011000101)
  ) CON2D_448(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[27][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111100001100111001010001111101)
)   op28(
    .i_pipeline_layer4(i_CORE_IP1[27]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*28-1:DATA_WIDTH*27])
);

/// CON2D_29///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001000011100110101101),
      .k2(32'b10111101110111100110001001011111),
      .k3(32'b10111101101000011111011101111011),
      .k4(32'b00111101100101001000101011011101),
      .k5(32'b10111001111110001111111001010100),
      .k6(32'b10111101110011100001100110111110),
      .k7(32'b10111101001010001101110001011111),
      .k8(32'b00111100100010001100001001111110),
      .k9(32'b10111100100101111111011010000001)
  ) CON2D_449(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111110000000101111010101010011),
      .k2(32'b10111101111000110111110000101110),
      .k3(32'b10111101000100010100011011000001),
      .k4(32'b10111101001001011101111110110011),
      .k5(32'b00111100110111111011110101111110),
      .k6(32'b10111101011111010110110000101111),
      .k7(32'b00111100001000101111110010101110),
      .k8(32'b10111100111011111101011000101110),
      .k9(32'b10111101111100000011011011011000)
  ) CON2D_450(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110011101011111010001100),
      .k2(32'b00111100000001100010111010111101),
      .k3(32'b00111101110010001100000001001011),
      .k4(32'b00111101101110010000100100111101),
      .k5(32'b10111101110111010110110000001000),
      .k6(32'b00111101101011110001100100100111),
      .k7(32'b10111011111001101011110111011100),
      .k8(32'b10111101011110100110110001010110),
      .k9(32'b00111101111000010001101010100000)
  ) CON2D_451(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010011011111100011001111),
      .k2(32'b00111100011110111001100010110010),
      .k3(32'b00111101111010001111001011010101),
      .k4(32'b10111101101110100010011101011101),
      .k5(32'b10111101011101001101101111000011),
      .k6(32'b10111101100011110001000100110000),
      .k7(32'b10111101110001001110001101110101),
      .k8(32'b00111101011111010011010001010110),
      .k9(32'b00111100100001001011011110000010)
  ) CON2D_452(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111010111011011110101100),
      .k2(32'b00111101100101100010001100011101),
      .k3(32'b00111101001001000100010011001100),
      .k4(32'b10111011001010000011110110100010),
      .k5(32'b00111100100001110000010110001001),
      .k6(32'b10111101101010101011011000100101),
      .k7(32'b00111101100110010101011111100001),
      .k8(32'b10111101000010010111010110011010),
      .k9(32'b10111110000011000111111100000000)
  ) CON2D_453(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000000001111101111100000),
      .k2(32'b00111100100101011001101111010010),
      .k3(32'b10111101010100111010111011111110),
      .k4(32'b00111100000000010111110010010110),
      .k5(32'b00111101110001011000000110101011),
      .k6(32'b00111100000100100001001010110010),
      .k7(32'b00111101000011101101101111011110),
      .k8(32'b00111100100110000010111011011001),
      .k9(32'b00111101101100001111111000011001)
  ) CON2D_454(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100000001011001011111111),
      .k2(32'b10111101101110011011001011101001),
      .k3(32'b10111101101011000001110110000000),
      .k4(32'b00111100111100110101100001110110),
      .k5(32'b00111100111001110111000010010110),
      .k6(32'b00111101000001110001100100000010),
      .k7(32'b00111100110001101010001001001011),
      .k8(32'b00111110000001011001111101110000),
      .k9(32'b10111011111100100001111101110000)
  ) CON2D_455(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110011111100100101101110),
      .k2(32'b10111101001111000111100011011011),
      .k3(32'b10111101111010010111111001111011),
      .k4(32'b10111101011010111010100000000001),
      .k5(32'b10111011111000010010000101101111),
      .k6(32'b10111101100100110010110011011001),
      .k7(32'b10111101010001010001110010100001),
      .k8(32'b00111100000111111010000100011000),
      .k9(32'b10111101111011101101011111111010)
  ) CON2D_456(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110000100110111011111000),
      .k2(32'b10111011110000000001100010011000),
      .k3(32'b00111011010000010101100110000101),
      .k4(32'b10111101001110110010100011111100),
      .k5(32'b10111100101101000010010100011100),
      .k6(32'b10111101100111010010100011011110),
      .k7(32'b10111101100100001000100111001011),
      .k8(32'b00111101110001000010110000011011),
      .k9(32'b00111101100001010010001011010001)
  ) CON2D_457(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111011111010011110100101110100),
      .k2(32'b10111101101000001110010101000011),
      .k3(32'b10111101100001001111000110100010),
      .k4(32'b10111101010001001010000000011011),
      .k5(32'b10111101000011001011010111001101),
      .k6(32'b00111101011101001101101111111001),
      .k7(32'b00111011011011001110111111011111),
      .k8(32'b00111101000110011001001101001010),
      .k9(32'b00111101001100101011000110101010)
  ) CON2D_458(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100111001011010111011101011),
      .k2(32'b10111101100111101101110010100000),
      .k3(32'b00111101010011000111100100101101),
      .k4(32'b10111101110001110000010001010000),
      .k5(32'b10111101100101100001000101110000),
      .k6(32'b10111011001001111101111111000001),
      .k7(32'b10111011000001101110010110100100),
      .k8(32'b10111101101000111001011110000110),
      .k9(32'b00111101111101011000010101000100)
  ) CON2D_459(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001011001100011111100),
      .k2(32'b10111101101100110011100101010011),
      .k3(32'b00111101111011001111001001000111),
      .k4(32'b00111101101001000100001100011100),
      .k5(32'b10111101101100111010011010110011),
      .k6(32'b10111101110111000101001110001011),
      .k7(32'b10111101110001101100110001101011),
      .k8(32'b10111101100000100000011100000001),
      .k9(32'b10111101011110000100010011110101)
  ) CON2D_460(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100100100101110111111000),
      .k2(32'b10111101011101100101110010010010),
      .k3(32'b10111101110011111100100001111000),
      .k4(32'b10111101000011100111111000100010),
      .k5(32'b00111101110100011110000011011111),
      .k6(32'b10111101100010101110101100010111),
      .k7(32'b10111100001100110001001101111100),
      .k8(32'b00111101110100101101011010100001),
      .k9(32'b00111100110110010011011001000110)
  ) CON2D_461(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111011000110101001100010),
      .k2(32'b10111101110101100000011000001100),
      .k3(32'b10111101101110100100110000111110),
      .k4(32'b10111100100100111101000110101011),
      .k5(32'b10111100110100000111111101110100),
      .k6(32'b00111101000000001110110110110101),
      .k7(32'b00111101100100010100001100111110),
      .k8(32'b00111100001001000111111010001111),
      .k9(32'b10111101011000011000111100111010)
  ) CON2D_462(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101111001001011000011011),
      .k2(32'b10111101101010000111001100011111),
      .k3(32'b00111011111110010000110111010001),
      .k4(32'b10111101110101111001010110110011),
      .k5(32'b00111101000011111100001101001101),
      .k6(32'b10111100011101001100111110111011),
      .k7(32'b10111100101100011110111011010100),
      .k8(32'b10111101000000010111100111000100),
      .k9(32'b00111101110011011010010011111111)
  ) CON2D_463(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100001011100010010011111),
      .k2(32'b10111101010010010101011010010000),
      .k3(32'b10111101100011110100110000100000),
      .k4(32'b00111101111101000000110101011101),
      .k5(32'b00111101001011001001110100010000),
      .k6(32'b10111101110010100111110010011101),
      .k7(32'b00111101001101100011001110111110),
      .k8(32'b10111101000001100101010100000011),
      .k9(32'b10111100101011101010100011001111)
  ) CON2D_464(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[28][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100010101010011001010100001)
)   op29(
    .i_pipeline_layer4(i_CORE_IP1[28]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*29-1:DATA_WIDTH*28])
);

/// CON2D_30///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101111001000110000110111001),
      .k2(32'b00111101101001011011100101011110),
      .k3(32'b00111100000010100010100010101111),
      .k4(32'b00111100010101011101110110000100),
      .k5(32'b00111100100100110101001111001110),
      .k6(32'b10111101110110010011011110011100),
      .k7(32'b10111011110011010010000100011010),
      .k8(32'b10111101010011111111111101100011),
      .k9(32'b10111100110010111011101101111000)
  ) CON2D_465(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111000100011000000101000),
      .k2(32'b10111100101000001001100101100001),
      .k3(32'b00111101010000111111100111001110),
      .k4(32'b00111101000100101010011011100011),
      .k5(32'b00111101100110100111000011111111),
      .k6(32'b10111100100100100000001100000110),
      .k7(32'b10111101011011011010110111101000),
      .k8(32'b10111101001110010010111001100010),
      .k9(32'b00111101101001101111000001100010)
  ) CON2D_466(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000011011010111010000100),
      .k2(32'b10111100111100110101100101100000),
      .k3(32'b00111101000000010101111001000111),
      .k4(32'b10111101100001101011101111110101),
      .k5(32'b00111101110010111011011000000010),
      .k6(32'b10111101101011110010110101000100),
      .k7(32'b10111101001001011111011000100011),
      .k8(32'b00111100011111011111011101011110),
      .k9(32'b00111101000110100000100001100111)
  ) CON2D_467(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100000110000010010000011),
      .k2(32'b10111100111111100100101000011101),
      .k3(32'b10111101101101000101110101011011),
      .k4(32'b10111101100110100000110100010011),
      .k5(32'b00111101000100010111000011100000),
      .k6(32'b00111101101011001110001011111011),
      .k7(32'b10111101110110100111001101100000),
      .k8(32'b00111101000101011010011101011111),
      .k9(32'b10111101100001001000001101001110)
  ) CON2D_468(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111011001111011011010100),
      .k2(32'b10111101001011101011111111100100),
      .k3(32'b00111101000110110111000110100000),
      .k4(32'b10111101010100101010010111110010),
      .k5(32'b10111101001001100110101001010000),
      .k6(32'b00111101110001001010011010011111),
      .k7(32'b00111101110000110101101011010110),
      .k8(32'b00111100111111011100001000001101),
      .k9(32'b10111101100110100101011010100100)
  ) CON2D_469(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110011101011000101001011),
      .k2(32'b10111101000000101100001111000111),
      .k3(32'b00111101111101101011101001000011),
      .k4(32'b10111101111101110110010010011101),
      .k5(32'b10111101001001101110000011111101),
      .k6(32'b00111010011001111010110000010010),
      .k7(32'b00111100101110011110010001101111),
      .k8(32'b00111101011001011011000001111111),
      .k9(32'b10111101000111100010010101001111)
  ) CON2D_470(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100111000000110011110),
      .k2(32'b00111101101100000111010010111110),
      .k3(32'b00111101110101111111101110111100),
      .k4(32'b10111101010010111001110100110000),
      .k5(32'b00111101000110101100111110011100),
      .k6(32'b00111101101001100101000001000110),
      .k7(32'b00111101100101101101011011100111),
      .k8(32'b00111100111110001001100101101100),
      .k9(32'b10111101100011111011000010000101)
  ) CON2D_471(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001100111111101011101111),
      .k2(32'b00111101011000001000010111001100),
      .k3(32'b00111100101011001111001000110010),
      .k4(32'b00111011101111010010100110101110),
      .k5(32'b10111101101001011111011001011001),
      .k6(32'b10111100101001000001011011010001),
      .k7(32'b00111101111011001110100111111001),
      .k8(32'b00111101100000111111000101110000),
      .k9(32'b00111101000100000111100010000001)
  ) CON2D_472(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010101001011111011000),
      .k2(32'b10111100011010000001010010001000),
      .k3(32'b00111101101111101100101000100010),
      .k4(32'b00111101001101001100111100011110),
      .k5(32'b00111100011000011011000111010011),
      .k6(32'b10111101011001010111010000000110),
      .k7(32'b10111101110010011101100011011000),
      .k8(32'b00111100100001110011111101111100),
      .k9(32'b10111101101111101010010000001000)
  ) CON2D_473(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101100001110011110001111),
      .k2(32'b00111100111011100110011101010111),
      .k3(32'b00111101110100110101001010110111),
      .k4(32'b00111101101011100110000011011010),
      .k5(32'b10111100111101100100000101111111),
      .k6(32'b10111101011001101011100011010011),
      .k7(32'b00111101101001100011001110011110),
      .k8(32'b00111101111100000011111000110101),
      .k9(32'b10111101001111010111011011011100)
  ) CON2D_474(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100011001000001111001001101),
      .k2(32'b00111101100100001101100110011011),
      .k3(32'b10111101100100101111011001101111),
      .k4(32'b00111100000010100010010100010111),
      .k5(32'b00111101010110011001100000011000),
      .k6(32'b00111101010000000001100011111111),
      .k7(32'b00111101010011011010100010110010),
      .k8(32'b10111101000000010110110100101010),
      .k9(32'b00111101101011110111001000011001)
  ) CON2D_475(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110011100111101001110100),
      .k2(32'b00111101101110111010000010011011),
      .k3(32'b10111100010010101001110111101001),
      .k4(32'b10111101001100001111111101011100),
      .k5(32'b00111110000010000011001111101001),
      .k6(32'b00111101101001001000110100101011),
      .k7(32'b10111101001100110000010001001101),
      .k8(32'b00111010111110100111111000100110),
      .k9(32'b00111101100101110100001000011010)
  ) CON2D_476(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001111110100101001010010),
      .k2(32'b10111101001010000011101111110111),
      .k3(32'b10111101011101100010000011110101),
      .k4(32'b10111101000110100110000110011100),
      .k5(32'b10111101001111010100101011110001),
      .k6(32'b10111011111011010100110011100110),
      .k7(32'b00111101010010001001000000110100),
      .k8(32'b00111101000110010111010111000101),
      .k9(32'b00111101100001110011010110010001)
  ) CON2D_477(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100111011110111110010010),
      .k2(32'b10111100101100001111000100000011),
      .k3(32'b10111100110000100010110000011010),
      .k4(32'b10111101000001100111001000000100),
      .k5(32'b00111011111110010001010010111110),
      .k6(32'b00111100111101101101011110111011),
      .k7(32'b10111101100000011011101110110000),
      .k8(32'b10111100111011101010101000010101),
      .k9(32'b00111100111111010011110101010011)
  ) CON2D_478(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100001110011000000011111),
      .k2(32'b10111100010101101001011101110101),
      .k3(32'b10111101000101000001001101000010),
      .k4(32'b10111101100110111000100101000000),
      .k5(32'b10111101100100011111110101110110),
      .k6(32'b10111010110111001010000111001111),
      .k7(32'b00111100110110000010011011100111),
      .k8(32'b10111101110110101110000110010101),
      .k9(32'b00111101101001100101000010011010)
  ) CON2D_479(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101100110110111101010110000),
      .k2(32'b00111101110010100110000011000110),
      .k3(32'b00111101111111011101011011100011),
      .k4(32'b00111101001100001010101010110001),
      .k5(32'b00111011101111100000111001010100),
      .k6(32'b10111101001010010111110011010100),
      .k7(32'b10111011111100000000001010010011),
      .k8(32'b10111101101101110000110000110000),
      .k9(32'b00111101111010000001110111000110)
  ) CON2D_480(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[29][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b00111100010101100010100101110010)
)   op30(
    .i_pipeline_layer4(i_CORE_IP1[29]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*30-1:DATA_WIDTH*29])
);

/// CON2D_31///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100101000011000010110111),
      .k2(32'b00111101010011111010100111010011),
      .k3(32'b00111101101001111010000000101011),
      .k4(32'b00111100000110101110100001100011),
      .k5(32'b00111101111011110000110010101001),
      .k6(32'b10111101100001000001100111000000),
      .k7(32'b00111101100010111100001001011101),
      .k8(32'b10111101100110010100011001001111),
      .k9(32'b00111100010000000100011010110101)
  ) CON2D_481(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000001111010101110010110),
      .k2(32'b00111101101100001011001100110101),
      .k3(32'b10111101100001101000100100000111),
      .k4(32'b10111101101011101001111011100000),
      .k5(32'b10111101100011001110000110100011),
      .k6(32'b00111101001011010100011111011001),
      .k7(32'b00111011110100011011110111111101),
      .k8(32'b10111101110111100111100101111010),
      .k9(32'b00111101110010100001101110101010)
  ) CON2D_482(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101001001111011000101111010),
      .k2(32'b00111101000001010111000111100100),
      .k3(32'b10111100110101010001000111000011),
      .k4(32'b00111101100110000000110001110101),
      .k5(32'b10111100111011010000011101111111),
      .k6(32'b10111101000001110010110010101010),
      .k7(32'b10111101100101111001010110101010),
      .k8(32'b10111100010110010001001011100110),
      .k9(32'b00111101011110111001000111111111)
  ) CON2D_483(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111101101001111001110100),
      .k2(32'b10111101101100110111000111010110),
      .k3(32'b10111101101101111100100011001110),
      .k4(32'b00111101010010111001011000100010),
      .k5(32'b00111100110110000010110010001000),
      .k6(32'b00111101100110010100010110100101),
      .k7(32'b00111101110110111110000011011001),
      .k8(32'b10111101110001110111000100001010),
      .k9(32'b10111101100000111010110100001110)
  ) CON2D_484(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101000100111100010011011110),
      .k2(32'b00111101101110011011101010110111),
      .k3(32'b00111101110111011000100001100011),
      .k4(32'b00111101001000101101000111100100),
      .k5(32'b00111101110001101111101000000001),
      .k6(32'b10111101001110101001010000001100),
      .k7(32'b00111101011011011100000010000100),
      .k8(32'b10111101100110110010101000000001),
      .k9(32'b00111101100111011011000101010010)
  ) CON2D_485(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100111110001100111000000101),
      .k2(32'b10111011000101001101111011111111),
      .k3(32'b00111101100010010000111000010101),
      .k4(32'b00111101110111001010101100011101),
      .k5(32'b00111101100001111111100001001011),
      .k6(32'b10111100001011000110110001010100),
      .k7(32'b10111101011010110111111101111101),
      .k8(32'b10111101110111110110000001010101),
      .k9(32'b00111101101101011011001101101010)
  ) CON2D_486(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101110010000010001000001101),
      .k2(32'b00111100011110001001111100110110),
      .k3(32'b10111011100111100001111001010011),
      .k4(32'b00111010100001110011101000100010),
      .k5(32'b00111101101101011101111100010101),
      .k6(32'b00111101101101111110010011011010),
      .k7(32'b10111101010010010111100000101110),
      .k8(32'b10111101101100100010111011100010),
      .k9(32'b10111101011010111100111111100001)
  ) CON2D_487(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101011001000000011000110110),
      .k2(32'b10111101010111101100010011110101),
      .k3(32'b10111100001100011111011001110111),
      .k4(32'b00111101011000001100000001100001),
      .k5(32'b00111101100000111011100110000110),
      .k6(32'b00111101001100110001000101111110),
      .k7(32'b00111101111100011011111000010101),
      .k8(32'b10111100111100010000011101010100),
      .k9(32'b00111101101110000101011110101011)
  ) CON2D_488(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101001000111110110101010011),
      .k2(32'b10111101110111100001010111110010),
      .k3(32'b00111101100001111001001101011111),
      .k4(32'b10111101111001110010000111001001),
      .k5(32'b00111101101111100111011000100011),
      .k6(32'b10111101110000100010100100010110),
      .k7(32'b00110111110010101011100000011011),
      .k8(32'b00111101101101001111011010111110),
      .k9(32'b10111100100010001010100110011111)
  ) CON2D_489(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111000011000110011111101),
      .k2(32'b10111101101111111011011100110111),
      .k3(32'b00111101001001100111111001100110),
      .k4(32'b10111101110000001000100000011100),
      .k5(32'b10111101101010001001111011100100),
      .k6(32'b10111101010101011001100011010011),
      .k7(32'b00111101110010100011110100111010),
      .k8(32'b00111101011001111001111111000010),
      .k9(32'b10111101101100110100111001000111)
  ) CON2D_490(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110001110100010101110101),
      .k2(32'b00111101101001000011101010111001),
      .k3(32'b10111010111100011111101100001100),
      .k4(32'b00111101101000111110111000111000),
      .k5(32'b00111101101001111101010111000101),
      .k6(32'b10111101101100111011001100101000),
      .k7(32'b10111101101000000000000100000100),
      .k8(32'b10111100100001101101010101000011),
      .k9(32'b00111101111010000110001001000111)
  ) CON2D_491(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101000011010101110011011101),
      .k2(32'b10111101010101010111001000111000),
      .k3(32'b10111101111010001011001100000100),
      .k4(32'b10111101101011010011000010111110),
      .k5(32'b10111101011011001111100101011101),
      .k6(32'b00111101100000010110010110100100),
      .k7(32'b00111101001001110111000000000100),
      .k8(32'b10111101101111000100111110001110),
      .k9(32'b10111101100110001001100001110001)
  ) CON2D_492(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101100011111000011011000100),
      .k2(32'b00111101101001110100000000001010),
      .k3(32'b00111100111010100111010111010010),
      .k4(32'b10111100001001010011110010000010),
      .k5(32'b10111101010011111011010100111101),
      .k6(32'b10111101010010100001100101011100),
      .k7(32'b10111101010110001010010010001000),
      .k8(32'b10111101110111100110101101000110),
      .k9(32'b00111100101101011010101010000010)
  ) CON2D_493(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111010101101000111000100101111),
      .k2(32'b10111100110001000110101011110000),
      .k3(32'b10111101000111001110101101100100),
      .k4(32'b10111101101000111010110110010001),
      .k5(32'b10111101001111000000001111010000),
      .k6(32'b10111101001001101010100101101001),
      .k7(32'b00111100101000000011110001001100),
      .k8(32'b00111101100100011110010011011001),
      .k9(32'b00111101100101001111010101111100)
  ) CON2D_494(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110010010110001101111100),
      .k2(32'b00111101100100111010011001100101),
      .k3(32'b00111101100101101100110001110101),
      .k4(32'b10111101001010011111111000111011),
      .k5(32'b00111011000110110111110000010100),
      .k6(32'b00111011101110100101011001111101),
      .k7(32'b10111101110111101010111101000101),
      .k8(32'b10111101001001100000100000100011),
      .k9(32'b00111100100001010001111001010000)
  ) CON2D_495(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010001011001100110110010),
      .k2(32'b00111100101011100111011001110101),
      .k3(32'b10111101111010100000011101111111),
      .k4(32'b10111011100011101110000000111100),
      .k5(32'b10111101101011111011101010001111),
      .k6(32'b00111101010101000010000011110111),
      .k7(32'b10111100010001010111100011111100),
      .k8(32'b10111101001100011010011010101001),
      .k9(32'b10111101111010000101010101011100)
  ) CON2D_496(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[30][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111100001011011001011001110001)
)   op31(
    .i_pipeline_layer4(i_CORE_IP1[30]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*31-1:DATA_WIDTH*30])
);

/// CON2D_32///////////////////
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100100111011011111101010100),
      .k2(32'b00111101111101011010101101001110),
      .k3(32'b00111101011001000011000000111110),
      .k4(32'b00111101101101101011100100101010),
      .k5(32'b10111100110111111011100100101011),
      .k6(32'b10111101110110011001011011101001),
      .k7(32'b00111101110100000111111001011101),
      .k8(32'b00111101111001100010000010001011),
      .k9(32'b10111101010110110010101101010001)
  ) CON2D_497(
      .i_data(i_data[DATA_WIDTH*1-1:DATA_WIDTH*0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*1-1:DATA_WIDTH*0])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101111000111111111100000000),
      .k2(32'b00111010100011101110011111100000),
      .k3(32'b10111101011011110100010001111011),
      .k4(32'b10111100101101111000101111111100),
      .k5(32'b10111101100001001100100001000100),
      .k6(32'b00111101101110011010011111001001),
      .k7(32'b00111100100000111111100110011010),
      .k8(32'b10111101000000000110010010111100),
      .k9(32'b10111011101111010110011011110000)
  ) CON2D_498(
      .i_data(i_data[DATA_WIDTH*2-1:DATA_WIDTH*1]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*2-1:DATA_WIDTH*1])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100110101011111001001001000),
      .k2(32'b00111101110011100110100100101101),
      .k3(32'b10111101101001101000101001010000),
      .k4(32'b10111101110001001010111100001000),
      .k5(32'b10111101111000101111101110010101),
      .k6(32'b10111101001010101110001011111101),
      .k7(32'b00111101001010001100100011011110),
      .k8(32'b00111101010011000001101010011000),
      .k9(32'b00111101110110001001111101010110)
  ) CON2D_499(
      .i_data(i_data[DATA_WIDTH*3-1:DATA_WIDTH*2]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*3-1:DATA_WIDTH*2])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111100011110101011111001101100),
      .k2(32'b00111101011001001010101110111010),
      .k3(32'b10111101010100100111101110000010),
      .k4(32'b10111101101100001011110101011010),
      .k5(32'b10111100011010000100011001011100),
      .k6(32'b00111101111011101110001010011110),
      .k7(32'b10111100111110000110011100100111),
      .k8(32'b00111011110100111100001110111111),
      .k9(32'b10111100010001101011010011111000)
  ) CON2D_500(
      .i_data(i_data[DATA_WIDTH*4-1:DATA_WIDTH*3]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*4-1:DATA_WIDTH*3])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110010101110001101001),
      .k2(32'b10111101100000010011100100111100),
      .k3(32'b00111101000100000011001000111100),
      .k4(32'b10111101110101100000100001101110),
      .k5(32'b10111101110100111000001010000001),
      .k6(32'b10111110000011010111010000110001),
      .k7(32'b10111101111111011100110100101110),
      .k8(32'b00111101110001111111010000110110),
      .k9(32'b10111101100100101110011010110110)
  ) CON2D_501(
      .i_data(i_data[DATA_WIDTH*5-1:DATA_WIDTH*4]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*5-1:DATA_WIDTH*4])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000000001000011100000101),
      .k2(32'b00111100101010001000100001111011),
      .k3(32'b00111101100000001011000101101000),
      .k4(32'b10111100101001101111111101110111),
      .k5(32'b00111100101010001001110100011111),
      .k6(32'b10111101000110001011011000011001),
      .k7(32'b10111101100110010000011010011110),
      .k8(32'b10111101101001101001110010100110),
      .k9(32'b00111101011001001110001101001101)
  ) CON2D_502(
      .i_data(i_data[DATA_WIDTH*6-1:DATA_WIDTH*5]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*6-1:DATA_WIDTH*5])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011111111100001010111110),
      .k2(32'b00111101110100010100011100110101),
      .k3(32'b00111101101010110100111101110001),
      .k4(32'b10111101100110100010111111010011),
      .k5(32'b10111101100101100101000001010110),
      .k6(32'b10111100100110111000110111001101),
      .k7(32'b10111101100111010001000000111000),
      .k8(32'b10111101010100100110101010110110),
      .k9(32'b10111100101000011101001001011010)
  ) CON2D_503(
      .i_data(i_data[DATA_WIDTH*7-1:DATA_WIDTH*6]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*7-1:DATA_WIDTH*6])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101110100111000110101010011),
      .k2(32'b00111101000110011010001110000101),
      .k3(32'b00111101111011101101101000000110),
      .k4(32'b10111100100101011101011010010100),
      .k5(32'b00111100101111110110001111111110),
      .k6(32'b00111101110111010100111010100100),
      .k7(32'b10111101101111110111010000000011),
      .k8(32'b10111011100001000000110011101101),
      .k9(32'b10111101011001111111100011110100)
  ) CON2D_504(
      .i_data(i_data[DATA_WIDTH*8-1:DATA_WIDTH*7]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*8-1:DATA_WIDTH*7])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111011001101101100001000110010),
      .k2(32'b00111101111011010011011001000101),
      .k3(32'b00111101100010000100001101011111),
      .k4(32'b00111011111001000100100111111111),
      .k5(32'b00111101100111000001000110001110),
      .k6(32'b00111011101000010010110110000100),
      .k7(32'b10111101100001010000001100001000),
      .k8(32'b10111101101000011011010101000101),
      .k9(32'b10111101100101100001001110111010)
  ) CON2D_505(
      .i_data(i_data[DATA_WIDTH*9-1:DATA_WIDTH*8]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*9-1:DATA_WIDTH*8])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101100001111011110100000),
      .k2(32'b00111101110001010110100000010000),
      .k3(32'b00111101001001010110010000110101),
      .k4(32'b00111101111010001001111001101011),
      .k5(32'b10111101000100001010110001110111),
      .k6(32'b10111101110110110100110011001110),
      .k7(32'b10111101001100111110000000001011),
      .k8(32'b00111101011100101101000000010011),
      .k9(32'b10111101110011001000101111011001)
  ) CON2D_506(
      .i_data(i_data[DATA_WIDTH*10-1:DATA_WIDTH*9]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*10-1:DATA_WIDTH*9])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111110000000001101001101011100),
      .k2(32'b10111100111010011111001011011111),
      .k3(32'b00111100001101101110100101100000),
      .k4(32'b10111101110001110000100011101100),
      .k5(32'b00111101110000111010000011101000),
      .k6(32'b00111101100111010100100010000011),
      .k7(32'b00111100010111000010100101111010),
      .k8(32'b00111101000111111010110111111011),
      .k9(32'b00111101011110010011110011001100)
  ) CON2D_507(
      .i_data(i_data[DATA_WIDTH*11-1:DATA_WIDTH*10]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*11-1:DATA_WIDTH*10])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111100100001010000110110100010),
      .k2(32'b10111101111000001011111101101001),
      .k3(32'b10111101011001010100101101001010),
      .k4(32'b10111100110100000100011101100110),
      .k5(32'b00111101101100111110011010111100),
      .k6(32'b00111100000101001000100101101100),
      .k7(32'b00111101101111010101100100111001),
      .k8(32'b00111101011100000100011111000001),
      .k9(32'b10111100001101111011011100011101)
  ) CON2D_508(
      .i_data(i_data[DATA_WIDTH*12-1:DATA_WIDTH*11]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*12-1:DATA_WIDTH*11])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101101100100000111000100111),
      .k2(32'b10111101011001010100001011110001),
      .k3(32'b00111001100100111001011011010100),
      .k4(32'b10111100001110000011110110011101),
      .k5(32'b00111101010101001110011010001100),
      .k6(32'b10111101101101110011000101100100),
      .k7(32'b00111100010101110010011010000111),
      .k8(32'b00111101000001000101010111110101),
      .k9(32'b00111101100111001100110000111110)
  ) CON2D_509(
      .i_data(i_data[DATA_WIDTH*13-1:DATA_WIDTH*12]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*13-1:DATA_WIDTH*12])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101101110101010001100110010),
      .k2(32'b10111101100001011010001011101011),
      .k3(32'b00111101100111111001000001100110),
      .k4(32'b00111101100110010100001100101100),
      .k5(32'b00111101100110000000011100011111),
      .k6(32'b10111101000110101101101010100111),
      .k7(32'b00111100010001111100111111101000),
      .k8(32'b00111101001111010100100110111100),
      .k9(32'b00111100100010101110100111101001)
  ) CON2D_510(
      .i_data(i_data[DATA_WIDTH*14-1:DATA_WIDTH*13]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*14-1:DATA_WIDTH*13])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b10111101011110101110111111001000),
      .k2(32'b10111101100101100101111011001010),
      .k3(32'b10111101001010001100011000110001),
      .k4(32'b00111101100001000101010001100110),
      .k5(32'b10111101101100000111000001100011),
      .k6(32'b00111101001000110000111010101001),
      .k7(32'b10111101101000001001001000010101),
      .k8(32'b00111101110001000011010110100010),
      .k9(32'b10111100000011111100111111011011)
  ) CON2D_511(
      .i_data(i_data[DATA_WIDTH*15-1:DATA_WIDTH*14]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*15-1:DATA_WIDTH*14])
  );

  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH),
      .k1(32'b00111101010111110100110010110000),
      .k2(32'b10111101001001110111100100111100),
      .k3(32'b10111101110111001101111001000000),
      .k4(32'b00111101101110101011111100100001),
      .k5(32'b10111101101110010101110000010010),
      .k6(32'b10111101000010000101010100111010),
      .k7(32'b10111101101010001001111111101010),
      .k8(32'b10111101111110010111110111111010),
      .k9(32'b10111010010100111111110000100001)
  ) CON2D_512(
      .i_data(i_data[DATA_WIDTH*16-1:DATA_WIDTH*15]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(padding_valid),
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .counter_col(counter_col),
      .counter_row(counter_row),
      .valid_pipeline2D(valid_pipeline2D),
      .o_data(i_CORE_IP1[31][DATA_WIDTH*16-1:DATA_WIDTH*15])
  );


pipeline_layer4#(
    .DATA_WIDTH(DATA_WIDTH),
    .bias(32'b10111010110010111001101101110011)
)   op32(
    .i_pipeline_layer4(i_CORE_IP1[31]), 
    .clk(clk),
    .rst(rst),
    .valid_in_bias(valid_in_bias),
    .valid_pipeline(valid_pipeline_bias),
    .o_data(o_data[DATA_WIDTH*32-1:DATA_WIDTH*31])
);

  control_layer5#(
      .WIDTH(WIDTH)
    )control( 
      .clk(clk), 
      .rst(rst),
      .valid_in(valid_in), 
      .padding_valid(padding_valid), 
      .counter_col(counter_col), 
      .counter_row(counter_row), 
      .valid_in_pipeline2D(valid_in_pipeline2D),
      .valid_pipeline2D(valid_pipeline2D),
      .valid_in_bias(valid_in_bias),
      .valid_pipeline_bias(valid_pipeline_bias),
      .valid_out(valid_out)
    );
endmodule
