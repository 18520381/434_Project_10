module layer15_1#(
  parameter DATA_WIDTH = 32
  )(
  input  [DATA_WIDTH*16-1:0] i_data,
  input         clk, rst, valid_in,
  output [DATA_WIDTH*2-1:0] o_data ,
  output valid_out
  );
  
  wire [4:0] valid_FC;

  FC_16#(
  .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110100111001101000100011101),
      .k2(32'b10111110100111011001111001000100),
      .k3(32'b10111110110100000000101110100000),
      .k4(32'b00111111000100000011000101010000),
      .k5(32'b00111101100000101001110010010000),
      .k6(32'b00111110010010111100000110010100),
      .k7(32'b10111110001110010000110100000011),
      .k8(32'b00111110011100001001000011001010),
      .k9(32'b00111110110100100001111011100100),
      .k10(32'b00111110111111110001111110100110),
      .k11(32'b00111110110011010101101111011101),
      .k12(32'b00111110101100110101100010010001),
      .k13(32'b10111110110010101010110111101000),
      .k14(32'b10111110000001101000000011000100),
      .k15(32'b00111010101010011110111010011000),
      .k16(32'b10111101111110110011010010111100),
      .bias(32'b00111100000101110011011110010001)
  ) FC1 (
      .i_data(i_data),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_FC),
      .o_data(o_data[DATA_WIDTH*1-1:DATA_WIDTH*0])  
  );

  FC_16#(
  .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110111000110100011111011000),
      .k2(32'b00111101101110100010111000001101),
      .k3(32'b00111110011011101011011001000011),
      .k4(32'b10111111000010100010010110010010),
      .k5(32'b00111110111111001100100011000101),
      .k6(32'b10111110100100101111100000010101),
      .k7(32'b10111110111111001101100101100100),
      .k8(32'b00111101100111111100110100011111),
      .k9(32'b00111111000010011101010010100100),
      .k10(32'b00111101011111100010011001100110),
      .k11(32'b10111110110100010111011110101100),
      .k12(32'b00111110111100011010010100101101),
      .k13(32'b10111110100010100101001000110101),
      .k14(32'b10111101101101000111111110100010),
      .k15(32'b00111101001001100101110011011000),
      .k16(32'b10111110110100101010100011100010),
      .bias(32'b10111100000101110011011110001101)
  ) FC2 (
      .i_data(i_data),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_FC),
      .o_data(o_data[DATA_WIDTH*2-1:DATA_WIDTH*1])  
  );

 control_FC_16 control1(
       .valid_in_FC(valid_in), 
       .clk(clk), 
       .rst(rst),
       .valid_out(valid_out),
       .valid_in_FC1(valid_FC)  
  );
endmodule

