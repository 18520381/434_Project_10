module layer1#(
    parameter DATA_WIDTH = 32,
    parameter WIDTH = 112,  
    parameter DEPTH = 12544 
)(
  input  [DATA_WIDTH*3-1:0] i_data,
  input              clk, rst, wr_req_FIFO_IN,
  output [DATA_WIDTH-1:0] o_data0, o_data1, o_data2, o_data3,
  output             valid_out            
);
  wire [DATA_WIDTH*3-1:0] o_fifo_in;
  wire empty_FIFO_IN, rd_req_FIFO_IN, valid_in_adder;
  wire [DATA_WIDTH-1:0]  o_CORE_IP1[63:0];
  wire [DATA_WIDTH-1:0]  o_CORE_IP2[63:0];
  wire [DATA_WIDTH-1:0]  o_CORE_IP3[63:0];
  wire [DATA_WIDTH-1:0]o_data4, o_data5, o_data6, o_data7, o_data8, o_data9, o_data10, o_data11, o_data12, o_data13, o_data14, o_data15, o_data16, o_data17, o_data18, o_data19, o_data20, o_data21, o_data22, o_data23, o_data24, o_data25, o_data26, o_data27, o_data28, o_data29, o_data30, o_data31, o_data32, o_data33, o_data34, o_data35, o_data36, o_data37, o_data38, o_data39, o_data40, o_data41, o_data42, o_data43, o_data44, o_data45, o_data46, o_data47, o_data48, o_data49, o_data50, o_data51, o_data52, o_data53, o_data54, o_data55, o_data56, o_data57, o_data58, o_data59, o_data60, o_data61, o_data62, o_data63;
  
  fifo #(
      .DATA_WIDTH(DATA_WIDTH),
      .DEPTH(DEPTH)
  ) FIFO_IN(
      .data_out(o_fifo_in),
      .empty(empty_FIFO_IN),
      .full(),
      .data_in(i_data),
      .wr_req(wr_req_FIFO_IN),
      .rd_req(rd_req_FIFO_IN),
      .rst(rst), 
      .clk(clk)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110110110111110001110010001),
      .k2(32'b00111111000011001110010110101011),
      .k3(32'b00111110111101011100010010010100),
      .k4(32'b00111110100011001010111010100011),
      .k5(32'b00111110101100010000010010110110),
      .k6(32'b00111110100111101111011011100000),
      .k7(32'b10111101011010110110001110111110),
      .k8(32'b10111101011100000010101100101010),
      .k9(32'b10111101010100000101111011010100)
  ) CON2D_1(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[0]),
      .valid_out(valid_in_adder),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101111110011011100010001),
      .k2(32'b00111110111000010101000101110011),
      .k3(32'b00111110110100010010110100100000),
      .k4(32'b00111101000111100110111110111100),
      .k5(32'b00111101001001100110110111110101),
      .k6(32'b00111101010011011010000011111111),
      .k7(32'b10111110100001100100010110010111),
      .k8(32'b10111110101010010100110110001001),
      .k9(32'b10111110100100100000100101010111)
  ) CON2D_2(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[0]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101011110110101010010111110),
      .k2(32'b10111101101001101010111000111111),
      .k3(32'b10111101100001010110101100001000),
      .k4(32'b10111110101111000000010010110011),
      .k5(32'b10111110111010000011000101010011),
      .k6(32'b10111110110011101000100001000110),
      .k7(32'b10111110101100110011111111100010),
      .k8(32'b10111110111110000101010111100001),
      .k9(32'b10111110110101100100011111000110)
  ) CON2D_3(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[0]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op0(
      .o_CORE_IP1(o_CORE_IP1[0]), 
      .o_CORE_IP2(o_CORE_IP2[0]), 
      .o_CORE_IP3(o_CORE_IP3[0]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data0), 
      .valid_out(valid_out)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111100000010110101001000),
      .k2(32'b00111100101010110000011100101001),
      .k3(32'b10111110001100001101011101100110),
      .k4(32'b00111110000101111110100100011011),
      .k5(32'b00111100111111100101101101000000),
      .k6(32'b10111110010000000001101010011011),
      .k7(32'b00111110000001000111001011010100),
      .k8(32'b00111101000000011100000110011001),
      .k9(32'b10111110001010011111110010011010)
  ) CON2D_4(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[1]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001001011111001110111111),
      .k2(32'b00111101010000011110100011100011),
      .k3(32'b10111110001011100111011011001100),
      .k4(32'b00111110010011110010011101010011),
      .k5(32'b00111101100001101100011110000010),
      .k6(32'b10111110001101011101010101010010),
      .k7(32'b00111110001011111011000010101110),
      .k8(32'b00111101011000000001011110110100),
      .k9(32'b10111110001010101010101010101111)
  ) CON2D_5(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[1]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000010101111001101011110),
      .k2(32'b00111101001010110110111110000001),
      .k3(32'b10111110000111100000111001010100),
      .k4(32'b00111110001001011001000110100110),
      .k5(32'b00111101001111010111100010000000),
      .k6(32'b10111110001100101001010111101000),
      .k7(32'b00111110000011100000101000011101),
      .k8(32'b00111101001011010101011101001101),
      .k9(32'b10111110001000001101000101100111)
  ) CON2D_6(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[1]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op1(
      .o_CORE_IP1(o_CORE_IP1[1]), 
      .o_CORE_IP2(o_CORE_IP2[1]), 
      .o_CORE_IP3(o_CORE_IP3[1]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data1), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101000010110101000100101100),
      .k2(32'b00111101110010100110011111111101),
      .k3(32'b00111101000110011101011000011110),
      .k4(32'b00111110001001010110111111110001),
      .k5(32'b00111110011101101000011101010000),
      .k6(32'b00111110001010101001011111111000),
      .k7(32'b00111100010100110110011100110010),
      .k8(32'b00111101100110111001000001001110),
      .k9(32'b00111100100000000000011000110000)
  ) CON2D_7(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[2]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111010110111111111010000101000),
      .k2(32'b00111101010100100111010111100000),
      .k3(32'b10111011101000101010000001110010),
      .k4(32'b00111110001000000010101100001111),
      .k5(32'b00111110011000011001100101010000),
      .k6(32'b00111110000110101101000100010011),
      .k7(32'b00111000011001000110011100101100),
      .k8(32'b00111101010001110110010001101101),
      .k9(32'b10111100000000101000011111101100)
  ) CON2D_8(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[2]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111011001111000100101000),
      .k2(32'b10111101110100000110100101000111),
      .k3(32'b10111110000011010101100111011010),
      .k4(32'b10111101101110000011000010100110),
      .k5(32'b10111101100010001011000011111110),
      .k6(32'b10111101111000001111100011011001),
      .k7(32'b10111110000000000101100100010100),
      .k8(32'b10111101111001011000100001000100),
      .k9(32'b10111110000110001011011001011000)
  ) CON2D_9(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[2]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op2(
      .o_CORE_IP1(o_CORE_IP1[2]), 
      .o_CORE_IP2(o_CORE_IP2[2]), 
      .o_CORE_IP3(o_CORE_IP3[2]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data2), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101101010101110001110010),
      .k2(32'b00111110110111111100001010110101),
      .k3(32'b00111110110100010100101100000010),
      .k4(32'b00111101110010000100101111011100),
      .k5(32'b00111101110001100001111100000100),
      .k6(32'b00111101110010110001100001000011),
      .k7(32'b10111010011111100111011101011000),
      .k8(32'b10111101010001010011100000011001),
      .k9(32'b10111100111000001001111101101110)
  ) CON2D_10(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[3]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100011101010110101000001),
      .k2(32'b00111110101001010011111110011011),
      .k3(32'b00111110101000010000010011111010),
      .k4(32'b10111110101110011000100000101011),
      .k5(32'b10111110110110010110110110011111),
      .k6(32'b10111110110010011111000110011000),
      .k7(32'b10111110110011100110110011000000),
      .k8(32'b10111111000000111111001001011110),
      .k9(32'b10111110111011111011101100101010)
  ) CON2D_11(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[3]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100110100111101110000010),
      .k2(32'b00111110101100111011100000010001),
      .k3(32'b00111110101100000110001110100110),
      .k4(32'b10111101001111001011110100010010),
      .k5(32'b10111101101101100010110110001011),
      .k6(32'b10111101011111010000001110000000),
      .k7(32'b10111110000101100101011110010111),
      .k8(32'b10111110011100001100000001000110),
      .k9(32'b10111110010001010111101010100000)
  ) CON2D_12(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[3]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op3(
      .o_CORE_IP1(o_CORE_IP1[3]), 
      .o_CORE_IP2(o_CORE_IP2[3]), 
      .o_CORE_IP3(o_CORE_IP3[3]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data3), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101101100010101001011001011),
      .k2(32'b10111101111000001111100111001101),
      .k3(32'b10111101101010000000000101001001),
      .k4(32'b10111110001111101111000111011010),
      .k5(32'b10111110011011111001110011001000),
      .k6(32'b10111110001110011100100000010101),
      .k7(32'b10111110011101010110001111000000),
      .k8(32'b10111110101011000111110011100000),
      .k9(32'b10111110100011100100100100101010)
  ) CON2D_13(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[4]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110010000110110110010010111),
      .k2(32'b00111110011101011100001000000001),
      .k3(32'b00111110100000000111111010001100),
      .k4(32'b00111110001101000101000001101001),
      .k5(32'b00111110010100101100111000100100),
      .k6(32'b00111110011110011010011001000111),
      .k7(32'b10111110000100001111111101011010),
      .k8(32'b10111110001101010111001010111001),
      .k9(32'b10111101111100001111111011101100)
  ) CON2D_14(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[4]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001011000111011011000110),
      .k2(32'b00111110011101000011111110111000),
      .k3(32'b00111110011011000010000111100000),
      .k4(32'b00111110000111011111011111110010),
      .k5(32'b00111110010101110110011101110001),
      .k6(32'b00111110011010011100000010101001),
      .k7(32'b10111101110100100100010000101001),
      .k8(32'b10111101111000000101101011001101),
      .k9(32'b10111101100010111000100010001111)
  ) CON2D_15(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[4]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op4(
      .o_CORE_IP1(o_CORE_IP1[4]), 
      .o_CORE_IP2(o_CORE_IP2[4]), 
      .o_CORE_IP3(o_CORE_IP3[4]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data4), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011010110011001000000010),
      .k2(32'b10111110010001001111111001111100),
      .k3(32'b10111101010001011100001000001101),
      .k4(32'b00111110100000001011100010000010),
      .k5(32'b10111110010101110110010110010000),
      .k6(32'b10111101100100101011100010101110),
      .k7(32'b00111110011001101000110110000110),
      .k8(32'b10111110010001010100001110001001),
      .k9(32'b10111101001110111101111111110001)
  ) CON2D_16(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[5]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011101010010011001001101),
      .k2(32'b10111110011001010000000111001101),
      .k3(32'b10111101101100000011101101110010),
      .k4(32'b00111110100010010000101110011001),
      .k5(32'b10111110011100011100001001100010),
      .k6(32'b10111101110100111000000001101001),
      .k7(32'b00111110100001010000100000001010),
      .k8(32'b10111110010010100010101000001100),
      .k9(32'b10111101011001100100111011111111)
  ) CON2D_17(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[5]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011011100000001101111111),
      .k2(32'b10111110001111111101111011000011),
      .k3(32'b10111101001100100000000100001001),
      .k4(32'b00111110011100101111001111111001),
      .k5(32'b10111110011000101111100110110101),
      .k6(32'b10111101101010001101010001100011),
      .k7(32'b00111110011000011011111100010100),
      .k8(32'b10111110010001101110111100101110),
      .k9(32'b10111101001111001011001001011111)
  ) CON2D_18(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[5]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op5(
      .o_CORE_IP1(o_CORE_IP1[5]), 
      .o_CORE_IP2(o_CORE_IP2[5]), 
      .o_CORE_IP3(o_CORE_IP3[5]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data5), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101100010001101111101101111),
      .k2(32'b00111101110010000111111001101011),
      .k3(32'b00111101100001100110001011101110),
      .k4(32'b00111110000101101100000010110101),
      .k5(32'b00111110010011011000111100010111),
      .k6(32'b00111110000111110011111111011001),
      .k7(32'b00111110000110111010110001001011),
      .k8(32'b00111110011010100111001110101010),
      .k9(32'b00111110001111000100011101010000)
  ) CON2D_19(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[6]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111001011000011000000010),
      .k2(32'b10111110000000001001100100100000),
      .k3(32'b10111110000101100111110100001011),
      .k4(32'b10111101010101111011111100010110),
      .k5(32'b10111101001100001010011001010100),
      .k6(32'b10111101100110110011010110100010),
      .k7(32'b00111101110010010010111001010101),
      .k8(32'b00111110000100001110001101010110),
      .k9(32'b00111101110101011100100010011000)
  ) CON2D_20(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[6]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001010101000001011011001),
      .k2(32'b10111110010101100010100001100100),
      .k3(32'b10111110010110001111111011101110),
      .k4(32'b10111110000111110101101111000100),
      .k5(32'b10111110001110000001001001010000),
      .k6(32'b10111110010001000001110011000011),
      .k7(32'b00111011111100100110110000110000),
      .k8(32'b00111100101001101000111111011100),
      .k9(32'b00111011100001010011010101010000)
  ) CON2D_21(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[6]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op6(
      .o_CORE_IP1(o_CORE_IP1[6]), 
      .o_CORE_IP2(o_CORE_IP2[6]), 
      .o_CORE_IP3(o_CORE_IP3[6]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data6), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001010010101001001101111),
      .k2(32'b00111101101000101000001100111110),
      .k3(32'b00111101111100011010100010001111),
      .k4(32'b10111110010110011011000101111110),
      .k5(32'b10111110011011101110001101111101),
      .k6(32'b10111110001011000001001010110011),
      .k7(32'b10111110010110100101010110110111),
      .k8(32'b10111110100100001001101000010110),
      .k9(32'b10111110011000101000111111110110)
  ) CON2D_22(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[7]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111011101100000000000010),
      .k2(32'b00111110010110011110101010101000),
      .k3(32'b00111110100000101011011010001100),
      .k4(32'b10111110000110001010000100110100),
      .k5(32'b10111101110110111011001010000100),
      .k6(32'b10111101000011111101000101001010),
      .k7(32'b10111110001111100010000011000100),
      .k8(32'b10111110010010111010001010001011),
      .k9(32'b10111110000000111010011110111100)
  ) CON2D_23(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[7]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110100110011000010100110),
      .k2(32'b00111110011100000101101010011101),
      .k3(32'b00111110100001101101110000101100),
      .k4(32'b00111101000111001010110001001110),
      .k5(32'b00111110000010010001000101101110),
      .k6(32'b00111110001111100101111010000001),
      .k7(32'b10111010110101100100101101110111),
      .k8(32'b00111101001011000001101011001011),
      .k9(32'b00111101101111110010110011010011)
  ) CON2D_24(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[7]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op7(
      .o_CORE_IP1(o_CORE_IP1[7]), 
      .o_CORE_IP2(o_CORE_IP2[7]), 
      .o_CORE_IP3(o_CORE_IP3[7]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data7), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000001010110010011101111),
      .k2(32'b10111110100011001110010000001101),
      .k3(32'b00111110001010000011100000110000),
      .k4(32'b00111101111001000001000011000011),
      .k5(32'b10111110100101100001101100110101),
      .k6(32'b00111110010010010100100100111101),
      .k7(32'b00111101110110011100111010111001),
      .k8(32'b10111110100100000011001101000001),
      .k9(32'b00111110001011111101111100000100)
  ) CON2D_25(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[8]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110001000101001001001100),
      .k2(32'b10111110101000110001011001101110),
      .k3(32'b00111110001011010101100111000000),
      .k4(32'b00111101100111100010001110101111),
      .k5(32'b10111110101010111100110011111011),
      .k6(32'b00111110010100010111110000111111),
      .k7(32'b00111101111010000100111010101100),
      .k8(32'b10111110100011111001111010001000),
      .k9(32'b00111110011000010010111100111000)
  ) CON2D_26(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[8]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000000010110010111011000),
      .k2(32'b10111110100011001001101010111101),
      .k3(32'b00111110001011010101100010001000),
      .k4(32'b00111101110010101101111100101111),
      .k5(32'b10111110100110011100101011111100),
      .k6(32'b00111110010001011101100011011001),
      .k7(32'b00111101110000010110000101010000),
      .k8(32'b10111110100100111001000000111010),
      .k9(32'b00111110001011010001011111011100)
  ) CON2D_27(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[8]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op8(
      .o_CORE_IP1(o_CORE_IP1[8]), 
      .o_CORE_IP2(o_CORE_IP2[8]), 
      .o_CORE_IP3(o_CORE_IP3[8]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data8), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101000001101100110100000000),
      .k2(32'b10111110000100011011111010100110),
      .k3(32'b10111110001000111001111100111111),
      .k4(32'b00111110000111001001111101010000),
      .k5(32'b10111100100000000010101101111001),
      .k6(32'b10111101011001101111000000110001),
      .k7(32'b00111110011011010011001011111001),
      .k8(32'b00111101110101110110100110111110),
      .k9(32'b00111101100010111001101000111001)
  ) CON2D_28(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[9]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101010101111011011011111001),
      .k2(32'b10111110100000001001011000101111),
      .k3(32'b10111110100011110011010001110100),
      .k4(32'b00111101110010001010010111001101),
      .k5(32'b10111101101111000010000011000100),
      .k6(32'b10111110000101000011011101010110),
      .k7(32'b00111110011110000110110000100100),
      .k8(32'b00111101110010011010110110001001),
      .k9(32'b00111101010000011011110011000010)
  ) CON2D_29(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[9]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100100000100100100101011111),
      .k2(32'b10111110001001001101000100010111),
      .k3(32'b10111110001110000010010011110001),
      .k4(32'b00111110000110001011101100101111),
      .k5(32'b10111100101010011110101011000100),
      .k6(32'b10111101100000001101001110101000),
      .k7(32'b00111110011010100100101011101000),
      .k8(32'b00111101110011111101010101111001),
      .k9(32'b00111101100000011011101000101001)
  ) CON2D_30(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[9]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op9(
      .o_CORE_IP1(o_CORE_IP1[9]), 
      .o_CORE_IP2(o_CORE_IP2[9]), 
      .o_CORE_IP3(o_CORE_IP3[9]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data9), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110001001110110010110000),
      .k2(32'b00111110001100010110001110110011),
      .k3(32'b00111110000101011010010011000111),
      .k4(32'b00111011011111000100110000001000),
      .k5(32'b00111100010001011010110100000001),
      .k6(32'b00111011010001111001011111101011),
      .k7(32'b10111110110001000001100000000101),
      .k8(32'b10111110111110100111011001010010),
      .k9(32'b10111110111010000000001011001101)
  ) CON2D_31(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[10]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111111000000000000110111111010),
      .k2(32'b00111111000110111100011110110011),
      .k3(32'b00111111000100001010001011110101),
      .k4(32'b00111110111110101100111111110010),
      .k5(32'b00111111000001110011111001011000),
      .k6(32'b00111111000000010110101001111110),
      .k7(32'b10111110101000000111101100110111),
      .k8(32'b10111110110100000011110111011110),
      .k9(32'b10111110101110110111111100001111)
  ) CON2D_32(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[10]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001111000101111100100000),
      .k2(32'b00111101111010000100000000011111),
      .k3(32'b00111101110010110111111111000011),
      .k4(32'b10111101001010100101100011011001),
      .k5(32'b10111101001100001001110101101011),
      .k6(32'b10111101000111000111100001111011),
      .k7(32'b10111110110001011111111000101110),
      .k8(32'b10111111000000000100011110001111),
      .k9(32'b10111110111010000100000000001101)
  ) CON2D_33(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[10]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op10(
      .o_CORE_IP1(o_CORE_IP1[10]), 
      .o_CORE_IP2(o_CORE_IP2[10]), 
      .o_CORE_IP3(o_CORE_IP3[10]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data10), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101101111001110000010100001),
      .k2(32'b00111101001010000001000011011000),
      .k3(32'b10111101101110010000111101010111),
      .k4(32'b10111110001000111010101111110011),
      .k5(32'b10111101010101100111010000010011),
      .k6(32'b10111110010000001101011010010101),
      .k7(32'b10111110011001100101100001010101),
      .k8(32'b10111110001010001010011000011001),
      .k9(32'b10111110100011010101111100011111)
  ) CON2D_34(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[11]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110101011100100000011011),
      .k2(32'b00111110100101101111000101011011),
      .k3(32'b00111110000010000111110001001101),
      .k4(32'b00111101101100110101011101010110),
      .k5(32'b00111110100000100100100000011000),
      .k6(32'b00111101101101010110011110101000),
      .k7(32'b10111110000110111111101010101010),
      .k8(32'b10111101001101111111010010100100),
      .k9(32'b10111110001110000011000101111010)
  ) CON2D_35(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[11]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001011001000010111110111),
      .k2(32'b00111110011110101110011100101110),
      .k3(32'b00111101101100111010010011101000),
      .k4(32'b00111101000111101101001100100111),
      .k5(32'b00111110011001000001010000100111),
      .k6(32'b00111101011101100110100111011111),
      .k7(32'b10111101111100001000001100111100),
      .k8(32'b00111100001100001000010011000101),
      .k9(32'b10111101111110100110011110001011)
  ) CON2D_36(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[11]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op11(
      .o_CORE_IP1(o_CORE_IP1[11]), 
      .o_CORE_IP2(o_CORE_IP2[11]), 
      .o_CORE_IP3(o_CORE_IP3[11]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data11), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000111111001110101000001),
      .k2(32'b00111110100101011100000111010100),
      .k3(32'b10111110011000000100100101110001),
      .k4(32'b10111110000100001001100011011010),
      .k5(32'b00111110101101110011100101010010),
      .k6(32'b10111110010000010001111100011011),
      .k7(32'b10111110001011111000000111100111),
      .k8(32'b00111110100110011111010010010110),
      .k9(32'b10111110010110011101110111011001)
  ) CON2D_37(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[12]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000100111100011100111110),
      .k2(32'b00111110101100100001000010100101),
      .k3(32'b10111110010010100010110010001011),
      .k4(32'b10111101110110010110000001001111),
      .k5(32'b00111110111000000001011001001000),
      .k6(32'b10111110000101000001011101101001),
      .k7(32'b10111110001000101100010100111101),
      .k8(32'b00111110101101010101100001010110),
      .k9(32'b10111110010001011011100100110010)
  ) CON2D_38(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[12]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000101110101101000111001),
      .k2(32'b00111110100111010110100010110001),
      .k3(32'b10111110010101101011110100001100),
      .k4(32'b10111101111111010111010001111101),
      .k5(32'b00111110110000100011111111111110),
      .k6(32'b10111110001100011110000000001100),
      .k7(32'b10111110001000100001001000000010),
      .k8(32'b00111110101000001011000110111100),
      .k9(32'b10111110010100110100100111010110)
  ) CON2D_39(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[12]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op12(
      .o_CORE_IP1(o_CORE_IP1[12]), 
      .o_CORE_IP2(o_CORE_IP2[12]), 
      .o_CORE_IP3(o_CORE_IP3[12]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data12), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101010101100011010100101011),
      .k2(32'b00111100100001011000000001011111),
      .k3(32'b10111110000000010011010000100101),
      .k4(32'b00111110010100000000100010111100),
      .k5(32'b00111110001101011110101111001100),
      .k6(32'b00111011100010101111100100001011),
      .k7(32'b00111110010011101011000010111011),
      .k8(32'b00111110010011010010000110110001),
      .k9(32'b00111101000111000011000001010110)
  ) CON2D_40(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[13]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111100011000011100011000000111),
      .k2(32'b10111101101000010000101110010101),
      .k3(32'b10111110011001111101010100100101),
      .k4(32'b00111110001100000000000010011010),
      .k5(32'b00111101111100101001001101010100),
      .k6(32'b10111101011101100110000000010011),
      .k7(32'b00111110010010101000001110001011),
      .k8(32'b00111110001100000101110000110010),
      .k9(32'b00111011010000111010110111011001)
  ) CON2D_41(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[13]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111001001001001001000110),
      .k2(32'b10111110001111111111010110001000),
      .k3(32'b10111110100111000011010000101101),
      .k4(32'b10111100101000010110010101000100),
      .k5(32'b10111101101101000100000011100110),
      .k6(32'b10111110011011011011101110011110),
      .k7(32'b00111101001011101010010111011101),
      .k8(32'b00111011011000100110111001011000),
      .k9(32'b10111110000001101110010011001011)
  ) CON2D_42(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[13]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op13(
      .o_CORE_IP1(o_CORE_IP1[13]), 
      .o_CORE_IP2(o_CORE_IP2[13]), 
      .o_CORE_IP3(o_CORE_IP3[13]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data13), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101101010100111101111101100),
      .k2(32'b10111110000000010001100100001110),
      .k3(32'b10111101110010111000010001111001),
      .k4(32'b10111101001100011001010001111101),
      .k5(32'b10111101010010101010010011111010),
      .k6(32'b10111100111111001010010000110101),
      .k7(32'b00111110011010101000001101111011),
      .k8(32'b00111110100111100110011111101110),
      .k9(32'b00111110100110001000010000010000)
  ) CON2D_43(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[14]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110110000110010110111010010),
      .k2(32'b10111110111010110000010100100110),
      .k3(32'b10111110110101011000111100011001),
      .k4(32'b10111110110011000110111111101001),
      .k5(32'b10111110110111111011001010111000),
      .k6(32'b10111110110011101111000011010011),
      .k7(32'b00111110001000101001000100000010),
      .k8(32'b00111110011001011111010111101010),
      .k9(32'b00111110011000110011111100111110)
  ) CON2D_44(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[14]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101011001001100011010100000),
      .k2(32'b10111101101011111011100110011101),
      .k3(32'b10111101011111001100010110100111),
      .k4(32'b00111100010000001011011000101100),
      .k5(32'b00111100101101011011000011101000),
      .k6(32'b00111101000100000001101000011111),
      .k7(32'b00111110100001101110100010110111),
      .k8(32'b00111110101101110101111010000010),
      .k9(32'b00111110101011100110111011010100)
  ) CON2D_45(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[14]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op14(
      .o_CORE_IP1(o_CORE_IP1[14]), 
      .o_CORE_IP2(o_CORE_IP2[14]), 
      .o_CORE_IP3(o_CORE_IP3[14]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data14), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001000010001000000000110),
      .k2(32'b10111110000111110100100101110110),
      .k3(32'b00111110001001000101100001000101),
      .k4(32'b00111101110011101000010100101001),
      .k5(32'b10111110011100011110001001100110),
      .k6(32'b00111101110100001001100100001000),
      .k7(32'b00111101111111011010001111001101),
      .k8(32'b10111110010011101011111111101101),
      .k9(32'b00111101110101001110000000011111)
  ) CON2D_46(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[15]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000011110000001010001100),
      .k2(32'b10111110010001011000111100100001),
      .k3(32'b00111110000110100111011101010111),
      .k4(32'b00111100111011011010101010101000),
      .k5(32'b10111110101010001110000010110010),
      .k6(32'b00111101000110011010101101111100),
      .k7(32'b00111101110101011010110001111011),
      .k8(32'b10111110011101010110000010110010),
      .k9(32'b00111101101111100010101000011010)
  ) CON2D_47(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[15]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000001001100001111001111),
      .k2(32'b10111110010000011010001101111111),
      .k3(32'b00111110000000010100100110100011),
      .k4(32'b00111101101101101010110000000100),
      .k5(32'b10111110100000001100010011011011),
      .k6(32'b00111101101011001011001111100111),
      .k7(32'b00111110000001001110001001111011),
      .k8(32'b10111110010010010111110011110001),
      .k9(32'b00111101110110000100011011110001)
  ) CON2D_48(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[15]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op15(
      .o_CORE_IP1(o_CORE_IP1[15]), 
      .o_CORE_IP2(o_CORE_IP2[15]), 
      .o_CORE_IP3(o_CORE_IP3[15]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data15), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100111011101000110000111000),
      .k2(32'b10111101010110011100101100111100),
      .k3(32'b00111110010000010011110001001010),
      .k4(32'b10111101001101110011011111001011),
      .k5(32'b10111101110000001101001100010111),
      .k6(32'b00111110011011010100100010111111),
      .k7(32'b10111101001011111100100100110110),
      .k8(32'b10111101110010101110111111001001),
      .k9(32'b00111110010110101011111111110101)
  ) CON2D_49(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[16]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101000001101111101100011110),
      .k2(32'b10111101110101101100010110100111),
      .k3(32'b00111110001110011001000010011000),
      .k4(32'b10111101111001011001011111110101),
      .k5(32'b10111110000110000011000101011101),
      .k6(32'b00111110011001110000100010100100),
      .k7(32'b10111101101001111011001111011100),
      .k8(32'b10111101111110111010100100001110),
      .k9(32'b00111110011100111000111011111111)
  ) CON2D_50(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[16]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101000100111100111010110100),
      .k2(32'b10111101011000000010101101010001),
      .k3(32'b00111110001101100001000110001001),
      .k4(32'b10111101000011110100111001110110),
      .k5(32'b10111101101110111000001001101110),
      .k6(32'b00111110011001101001011000010001),
      .k7(32'b10111101000100000110000111100001),
      .k8(32'b10111101110001001100111010110000),
      .k9(32'b00111110010101010111011111010000)
  ) CON2D_51(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[16]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op16(
      .o_CORE_IP1(o_CORE_IP1[16]), 
      .o_CORE_IP2(o_CORE_IP2[16]), 
      .o_CORE_IP3(o_CORE_IP3[16]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data16), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101010100001010111100111000),
      .k2(32'b00111110001110011010010111110111),
      .k3(32'b00111101101111110111000000000110),
      .k4(32'b00111101100100011010110111011101),
      .k5(32'b00111110010001001111001111101001),
      .k6(32'b00111101110010100100011111011111),
      .k7(32'b10111101101010100011111110101100),
      .k8(32'b10111010010001011100100110101110),
      .k9(32'b10111101100101010011010100001010)
  ) CON2D_52(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[17]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101101010111000000111010100),
      .k2(32'b00111110010010110010100001010000),
      .k3(32'b00111101111000010110011010001000),
      .k4(32'b00111101110101001101001110111001),
      .k5(32'b00111110010100110100111011101100),
      .k6(32'b00111101111001110000101111001011),
      .k7(32'b10111101110001101111110100010000),
      .k8(32'b10111101000011110101110111011001),
      .k9(32'b10111101110110101100001110011101)
  ) CON2D_53(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[17]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101101111101111111111011111),
      .k2(32'b10111100110100001010001000001000),
      .k3(32'b10111101101101111000001100010101),
      .k4(32'b10111110000101001100100000101010),
      .k5(32'b10111101101111100111101100011010),
      .k6(32'b10111110001001001100111011110011),
      .k7(32'b10111110001110111110001110000000),
      .k8(32'b10111110001001011100011110010110),
      .k9(32'b10111110010111000000111001010100)
  ) CON2D_54(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[17]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op17(
      .o_CORE_IP1(o_CORE_IP1[17]), 
      .o_CORE_IP2(o_CORE_IP2[17]), 
      .o_CORE_IP3(o_CORE_IP3[17]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data17), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110010000110010000110000000),
      .k2(32'b10111110010101001011010001011110),
      .k3(32'b00111101100110011000101110100110),
      .k4(32'b00111110010011100110010001011011),
      .k5(32'b10111110010111111001100101100011),
      .k6(32'b00111101101000000011101100010001),
      .k7(32'b00111110010001011011110100000100),
      .k8(32'b10111110010011001001010011111011),
      .k9(32'b00111101101011111001011111011011)
  ) CON2D_55(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[18]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001010101010110100101000),
      .k2(32'b10111110100001000010110110101111),
      .k3(32'b00111101001010110101111100001010),
      .k4(32'b00111101111001001110111000100001),
      .k5(32'b10111110101010111011111100001010),
      .k6(32'b10111100101000011110111000001111),
      .k7(32'b00111110000101110000000011000011),
      .k8(32'b10111110100010100011111001011111),
      .k9(32'b00111101000001111111000111001001)
  ) CON2D_56(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[18]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110010010111101011111100100),
      .k2(32'b10111110010010000000001101001110),
      .k3(32'b00111101101110010011110011111110),
      .k4(32'b00111110010110000101001110101001),
      .k5(32'b10111110010100000001010101100001),
      .k6(32'b00111101110000111100011111110011),
      .k7(32'b00111110010000110101000101111000),
      .k8(32'b10111110010010001100101111010010),
      .k9(32'b00111101101110111111010011101000)
  ) CON2D_57(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[18]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op18(
      .o_CORE_IP1(o_CORE_IP1[18]), 
      .o_CORE_IP2(o_CORE_IP2[18]), 
      .o_CORE_IP3(o_CORE_IP3[18]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data18), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101001100110001011000100100),
      .k2(32'b10111110000011100100011111101001),
      .k3(32'b00111110000000010101101100101110),
      .k4(32'b10111101101011011000000111010101),
      .k5(32'b10111110000101011101110111101011),
      .k6(32'b00111110010001100011111010011111),
      .k7(32'b10111101100000001001000011110000),
      .k8(32'b10111101111110110011110010010010),
      .k9(32'b00111110001110100010000000011011)
  ) CON2D_58(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[19]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101110101010101000111110001),
      .k2(32'b10111110010000111111001011011100),
      .k3(32'b00111110000000101100100011000101),
      .k4(32'b10111110000111111000011101001111),
      .k5(32'b10111110010101000000010011000101),
      .k6(32'b00111110010000101011001001111101),
      .k7(32'b10111101110011111101000111100111),
      .k8(32'b10111110000101110000011101100111),
      .k9(32'b00111110010110000110000001101111)
  ) CON2D_59(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[19]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101010000010000100011111101),
      .k2(32'b10111110000101001110101011111111),
      .k3(32'b00111101111011010101011001111010),
      .k4(32'b10111101101110010111000010111000),
      .k5(32'b10111110000111010110000010000001),
      .k6(32'b00111110001110110001110111011000),
      .k7(32'b10111101100100011110011001100100),
      .k8(32'b10111110000001100001110111111011),
      .k9(32'b00111110001011100101000010001111)
  ) CON2D_60(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[19]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op19(
      .o_CORE_IP1(o_CORE_IP1[19]), 
      .o_CORE_IP2(o_CORE_IP2[19]), 
      .o_CORE_IP3(o_CORE_IP3[19]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data19), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101110010011111001000010),
      .k2(32'b00111110100000101100001010011110),
      .k3(32'b00111110011101000011100100100010),
      .k4(32'b00111110100011010001101111110101),
      .k5(32'b00111101111101101101111111011011),
      .k6(32'b00111101110011011111011111010001),
      .k7(32'b00111110000010100011011110010010),
      .k8(32'b10111100111101110110010011111100),
      .k9(32'b10111100110100100110011111110000)
  ) CON2D_61(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[20]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100111011111001100111011),
      .k2(32'b00111110001000001000101001101111),
      .k3(32'b00111110000100001111100001110010),
      .k4(32'b00111101101110010110110111010001),
      .k5(32'b10111101111100011001010001100100),
      .k6(32'b10111110000001100011111111101011),
      .k7(32'b10111100110100011011101000010010),
      .k8(32'b10111110011110010111011001010011),
      .k9(32'b10111110011011110011111011000100)
  ) CON2D_62(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[20]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000011111110111101111110),
      .k2(32'b10111100101001001100001111000100),
      .k3(32'b10111011101110011100100101100001),
      .k4(32'b10111101100111000110100010011011),
      .k5(32'b10111110100101101001011001001110),
      .k6(32'b10111110100011100100110010110010),
      .k7(32'b10111110000100010000011111001100),
      .k8(32'b10111110101110101011001100000100),
      .k9(32'b10111110101010001011001010110011)
  ) CON2D_63(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[20]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op20(
      .o_CORE_IP1(o_CORE_IP1[20]), 
      .o_CORE_IP2(o_CORE_IP2[20]), 
      .o_CORE_IP3(o_CORE_IP3[20]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data20), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011101001100001111110011),
      .k2(32'b00111110101101100110111011101000),
      .k3(32'b00111110101101100100000111101111),
      .k4(32'b00111101101110000111011000010110),
      .k5(32'b00111110000101110111010101110000),
      .k6(32'b00111110001110101010110011001110),
      .k7(32'b10111010001110101000001011000101),
      .k8(32'b10111100001100101111010101111110),
      .k9(32'b00111101000011111000011111010110)
  ) CON2D_64(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[21]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100111101010011111111001),
      .k2(32'b00111110110000101000011100010111),
      .k3(32'b00111110110010111011011111100010),
      .k4(32'b10111101100110111101101100110001),
      .k5(32'b10111101101011010010010000001001),
      .k6(32'b10111100110011110010001101100010),
      .k7(32'b10111110010100100111111101000111),
      .k8(32'b10111110100100100101110110001100),
      .k9(32'b10111110010111100010000101100110)
  ) CON2D_65(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[21]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101100001001001010001101011),
      .k2(32'b00111101011010100010100111010101),
      .k3(32'b00111101101100010001011100000101),
      .k4(32'b10111110100000101110110001000110),
      .k5(32'b10111110101011111000010111001100),
      .k6(32'b10111110100011101111011110001000),
      .k7(32'b10111110100000000000011110100000),
      .k8(32'b10111110110010101010111100010101),
      .k9(32'b10111110101010011000010101111000)
  ) CON2D_66(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[21]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op21(
      .o_CORE_IP1(o_CORE_IP1[21]), 
      .o_CORE_IP2(o_CORE_IP2[21]), 
      .o_CORE_IP3(o_CORE_IP3[21]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data21), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001010101010110000001011),
      .k2(32'b00111010100110110101000101010100),
      .k3(32'b10111101111101101011010001110110),
      .k4(32'b00111110001101110110010001000001),
      .k5(32'b10111100100111000110111010101000),
      .k6(32'b10111110001001111010011010000111),
      .k7(32'b00111110001001000110001100001110),
      .k8(32'b10111100000111001110111000010001),
      .k9(32'b10111110000010010010100010111110)
  ) CON2D_67(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[22]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001011110001010011011100),
      .k2(32'b10111100110101001000010000010101),
      .k3(32'b10111110001011110000000011001000),
      .k4(32'b00111110001101111010011100110011),
      .k5(32'b10111101010100110111010110011001),
      .k6(32'b10111110011000001001100000000000),
      .k7(32'b00111110010001000000100110010101),
      .k8(32'b10111100001010101011111001100010),
      .k9(32'b10111110001000010000111001011011)
  ) CON2D_68(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[22]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001011001100010011110110),
      .k2(32'b00111010110001011111101100000100),
      .k3(32'b10111101111111100000110101110010),
      .k4(32'b00111110001011100101010110000100),
      .k5(32'b10111100111110001100110010011110),
      .k6(32'b10111110001101100010111001110100),
      .k7(32'b00111110001011001101101101111110),
      .k8(32'b10111011011110000011011111011100),
      .k9(32'b10111110000001011110101110010101)
  ) CON2D_69(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[22]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op22(
      .o_CORE_IP1(o_CORE_IP1[22]), 
      .o_CORE_IP2(o_CORE_IP2[22]), 
      .o_CORE_IP3(o_CORE_IP3[22]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data22), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001110001100110001110110),
      .k2(32'b10111110111110010101101110110111),
      .k3(32'b10111110100111011101111010000011),
      .k4(32'b10111101101000111010001111110011),
      .k5(32'b10111110110000000110100110111001),
      .k6(32'b10111110010100001000000111110110),
      .k7(32'b00111110001111001110110000110111),
      .k8(32'b10111101010001010011000100001100),
      .k9(32'b00111101110110110100000011101001)
  ) CON2D_70(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[23]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111100000001111000100101),
      .k2(32'b10111110110100011010101111000000),
      .k3(32'b10111110011100111001110101011111),
      .k4(32'b10111001101101110111100101101110),
      .k5(32'b10111110100011011101001010011000),
      .k6(32'b10111101111011111111100111100101),
      .k7(32'b00111110100011100001100110010101),
      .k8(32'b00111101100000001101101000101100),
      .k9(32'b00111110010100001000001111001000)
  ) CON2D_71(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[23]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001110011101011111101001),
      .k2(32'b10111101001100001100010101001011),
      .k3(32'b00111101110111100001110111011110),
      .k4(32'b00111110101011100010101101110110),
      .k5(32'b00111110000001011000011000100111),
      .k6(32'b00111110100010000110101101100111),
      .k7(32'b00111110110011110100011001010001),
      .k8(32'b00111110011110011001100001110011),
      .k9(32'b00111110101111001101010100000001)
  ) CON2D_72(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[23]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op23(
      .o_CORE_IP1(o_CORE_IP1[23]), 
      .o_CORE_IP2(o_CORE_IP2[23]), 
      .o_CORE_IP3(o_CORE_IP3[23]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data23), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001101000110101111100100),
      .k2(32'b00111101111011000011011001001001),
      .k3(32'b10111100101010101010101111111001),
      .k4(32'b00111101100110001001110001001100),
      .k5(32'b00111110000101101100100100110110),
      .k6(32'b10111010000001111111100010000011),
      .k7(32'b00111101001001001110001001011001),
      .k8(32'b00111101111010101100100001011011),
      .k9(32'b10111100101100111100011010000001)
  ) CON2D_73(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[24]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100000111100101001011101110),
      .k2(32'b00111101100010010011111011010100),
      .k3(32'b10111101100100101000100011100100),
      .k4(32'b00111100111000001110101111010000),
      .k5(32'b00111101101011100010100110000101),
      .k6(32'b10111101100000111110001000011000),
      .k7(32'b00111100011110010001011111110000),
      .k8(32'b00111101100110110101101010011111),
      .k9(32'b10111101100000010101000000111111)
  ) CON2D_74(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[24]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101001111000001100010100100),
      .k2(32'b10111011001000011100010000011110),
      .k3(32'b10111101111110100110111101111010),
      .k4(32'b10111101011100010010110111000010),
      .k5(32'b10111100100010110000010000000010),
      .k6(32'b10111110000101011110001001011101),
      .k7(32'b10111101001111000110000110110101),
      .k8(32'b00111001101110000110011000100001),
      .k9(32'b10111101111101010001110010011100)
  ) CON2D_75(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[24]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op24(
      .o_CORE_IP1(o_CORE_IP1[24]), 
      .o_CORE_IP2(o_CORE_IP2[24]), 
      .o_CORE_IP3(o_CORE_IP3[24]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data24), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110001000111011000011000),
      .k2(32'b00111101111011100101100001010011),
      .k3(32'b10111110001000101000100100100111),
      .k4(32'b00111101111110101000011001101010),
      .k5(32'b00111110000011001010101000100100),
      .k6(32'b10111110001010110101001010001011),
      .k7(32'b00111101101000101001000111101111),
      .k8(32'b00111101110101111000101100110110),
      .k9(32'b10111110001100011111100000011100)
  ) CON2D_76(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[25]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111111110101100001101101),
      .k2(32'b00111110000011101100101100011011),
      .k3(32'b10111110001001110001101110011001),
      .k4(32'b00111110000111000111001111011001),
      .k5(32'b00111110001001010010000001111101),
      .k6(32'b10111110001100001010011011001001),
      .k7(32'b00111101111011000010111000000000),
      .k8(32'b00111110000010001101011101111101),
      .k9(32'b10111110001100011000101101010100)
  ) CON2D_77(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[25]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110100000101110101100010),
      .k2(32'b00111110000000010110010011111010),
      .k3(32'b10111110000111000001000010010001),
      .k4(32'b00111110000001001011111110100111),
      .k5(32'b00111110000101101110100101010111),
      .k6(32'b10111110001001001111011101010101),
      .k7(32'b00111101101011101111111110001001),
      .k8(32'b00111101111001011111110100001111),
      .k9(32'b10111110001011101100000000011101)
  ) CON2D_78(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[25]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op25(
      .o_CORE_IP1(o_CORE_IP1[25]), 
      .o_CORE_IP2(o_CORE_IP2[25]), 
      .o_CORE_IP3(o_CORE_IP3[25]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data25), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101001100110111001101111100),
      .k2(32'b10111101100111011110000010001011),
      .k3(32'b10111101100100100110101110100100),
      .k4(32'b00111110001111100010001101011010),
      .k5(32'b00111110011101110000101110100101),
      .k6(32'b00111110011010010110101111000010),
      .k7(32'b00111110100010110100110101001001),
      .k8(32'b00111110110100010011011111111010),
      .k9(32'b00111110101111111100100011000000)
  ) CON2D_79(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[26]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110110010000011010100010101),
      .k2(32'b10111110111111010111010010110100),
      .k3(32'b10111110111100000100111101101001),
      .k4(32'b10111101110101010110110110101101),
      .k5(32'b10111101110111111010101101010111),
      .k6(32'b10111101110011100011000010011010),
      .k7(32'b00111110011111101111111001010000),
      .k8(32'b00111110101100001110100011010111),
      .k9(32'b00111110101001100100110100111101)
  ) CON2D_80(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[26]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100100100100000010101100),
      .k2(32'b10111110110101001101100100010101),
      .k3(32'b10111110110001101010111011110101),
      .k4(32'b10111101101101000111110011011100),
      .k5(32'b10111110000001001010111000000010),
      .k6(32'b10111101111011000011111000010110),
      .k7(32'b00111110001100100110010100010010),
      .k8(32'b00111110011011011011111111101101),
      .k9(32'b00111110011000101100001111001111)
  ) CON2D_81(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[26]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op26(
      .o_CORE_IP1(o_CORE_IP1[26]), 
      .o_CORE_IP2(o_CORE_IP2[26]), 
      .o_CORE_IP3(o_CORE_IP3[26]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data26), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110010000010000000111010010),
      .k2(32'b00111101110101000101100111011100),
      .k3(32'b10111101010011101001010001110000),
      .k4(32'b10111110001111010100000010000111),
      .k5(32'b00111110000100111001100000110101),
      .k6(32'b10111011101000000000110100111111),
      .k7(32'b10111110010001100000101000010010),
      .k8(32'b00111101101010110100101001010101),
      .k9(32'b10111101100001011011110000011001)
  ) CON2D_82(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[27]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001101100011001010011000),
      .k2(32'b00111110001100100101100011111001),
      .k3(32'b00111100110111110111100110010101),
      .k4(32'b10111110000001000000100111101011),
      .k5(32'b00111110100001110110110010110100),
      .k6(32'b00111101111110011101100000000100),
      .k7(32'b10111110001111100101100100000110),
      .k8(32'b00111110000101111011111111110001),
      .k9(32'b00111011111010001111101100000010)
  ) CON2D_83(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[27]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001110110101000011010111),
      .k2(32'b00111110000011110011100110101001),
      .k3(32'b10111011101101011101001111110011),
      .k4(32'b10111110001011100100001101001000),
      .k5(32'b00111110010000110001110101111110),
      .k6(32'b00111101010100000111001010000110),
      .k7(32'b10111110010000111110110010101110),
      .k8(32'b00111101111010000001110010100111),
      .k9(32'b10111100110110000101100100010011)
  ) CON2D_84(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[27]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op27(
      .o_CORE_IP1(o_CORE_IP1[27]), 
      .o_CORE_IP2(o_CORE_IP2[27]), 
      .o_CORE_IP3(o_CORE_IP3[27]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data27), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101001101000011010000100000),
      .k2(32'b10111101100100110010100111000100),
      .k3(32'b10111101000010101001101100111001),
      .k4(32'b10111110101100010010000111111100),
      .k5(32'b10111110110110000100111010101110),
      .k6(32'b10111110101111011001000100001100),
      .k7(32'b10111101100010101000010010010011),
      .k8(32'b10111101110101000000001110011100),
      .k9(32'b10111101100011000111100010001111)
  ) CON2D_85(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[28]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101000101110000110011110110),
      .k2(32'b10111100101110100101111010101001),
      .k3(32'b10111010111101011111111000001100),
      .k4(32'b10111110110111011010010101101000),
      .k5(32'b10111110111011100001110000110001),
      .k6(32'b10111110110111001000110101100010),
      .k7(32'b10111101101000001101000011110100),
      .k8(32'b10111101100100110110100111100111),
      .k9(32'b10111101011000101101001000001101)
  ) CON2D_86(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[28]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100011111101000010011101),
      .k2(32'b00111110110001100100101100001100),
      .k3(32'b00111110101111001101001110010000),
      .k4(32'b00111110010100011110000000010101),
      .k5(32'b00111110100100011111000000001000),
      .k6(32'b00111110100011000100001001100010),
      .k7(32'b00111110011101101000010011101101),
      .k8(32'b00111110101011011011001111001110),
      .k9(32'b00111110101000100011011101110001)
  ) CON2D_87(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[28]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op28(
      .o_CORE_IP1(o_CORE_IP1[28]), 
      .o_CORE_IP2(o_CORE_IP2[28]), 
      .o_CORE_IP3(o_CORE_IP3[28]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data28), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110010000100110100100110101),
      .k2(32'b10111011011111101001011110100100),
      .k3(32'b00111110011000001101011011101101),
      .k4(32'b10111110010001100111111011100001),
      .k5(32'b10111100011010001101101010101101),
      .k6(32'b00111110011010011010100101000010),
      .k7(32'b10111110001000101111010001111010),
      .k8(32'b10111101100001101111101000101011),
      .k9(32'b00111101110011111000011010000000)
  ) CON2D_88(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[29]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001101001001000110101011),
      .k2(32'b00111100101110011110110010101010),
      .k3(32'b00111110100010101011001010100000),
      .k4(32'b10111110001101101010010010001010),
      .k5(32'b00111100010001110000110101100111),
      .k6(32'b00111110100011101100110001111110),
      .k7(32'b10111110001111001111110010100101),
      .k8(32'b10111101101011001000011010010110),
      .k9(32'b00111101110101111110100010011010)
  ) CON2D_89(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[29]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001001000101110000010001),
      .k2(32'b10111100111011011100011101111111),
      .k3(32'b00111110000101001010100011110100),
      .k4(32'b10111110001011101111110100001010),
      .k5(32'b10111101010000110100001111111011),
      .k6(32'b00111110000100110000010010000111),
      .k7(32'b10111101111111101101010011111011),
      .k8(32'b10111101101000111100000111100100),
      .k9(32'b00111101000101000001011100000111)
  ) CON2D_90(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[29]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op29(
      .o_CORE_IP1(o_CORE_IP1[29]), 
      .o_CORE_IP2(o_CORE_IP2[29]), 
      .o_CORE_IP3(o_CORE_IP3[29]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data29), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110011011110111101110010010),
      .k2(32'b10111110100001101110101010001111),
      .k3(32'b10111110100101011000100111000000),
      .k4(32'b10111101110111110111110111101110),
      .k5(32'b10111101110010100111010101110011),
      .k6(32'b10111110000110100001110101101101),
      .k7(32'b10111101001001010011010100110100),
      .k8(32'b00111011001011110001001110100110),
      .k9(32'b10111101010011011011011011100111)
  ) CON2D_91(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[30]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001010111101011001110001),
      .k2(32'b10111110001010011010011111110010),
      .k3(32'b10111110010111001000000011011111),
      .k4(32'b00111110001011011100000001010000),
      .k5(32'b00111110011000101011001000110011),
      .k6(32'b00111110000011111011011010111000),
      .k7(32'b00111110001110000110110010111101),
      .k8(32'b00111110100001011110010100011001),
      .k9(32'b00111110001101111110110000001000)
  ) CON2D_92(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[30]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101110010011011111001100101),
      .k2(32'b10111101100100111010011101101110),
      .k3(32'b10111101111111000010101000100011),
      .k4(32'b00111110000001101000111101101111),
      .k5(32'b00111110010011110100100001100000),
      .k6(32'b00111101111110011110110110110001),
      .k7(32'b00111101111101011000000100010100),
      .k8(32'b00111110010111001001000100111001),
      .k9(32'b00111110000011001001010011100100)
  ) CON2D_93(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[30]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op30(
      .o_CORE_IP1(o_CORE_IP1[30]), 
      .o_CORE_IP2(o_CORE_IP2[30]), 
      .o_CORE_IP3(o_CORE_IP3[30]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data30), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000000110111001011000001),
      .k2(32'b00111101111111101110101111111011),
      .k3(32'b00111110000110001000001011110011),
      .k4(32'b00111101111000101010001010010001),
      .k5(32'b00111101111011101111110001001001),
      .k6(32'b00111110000100010001111010001000),
      .k7(32'b00111110001000111001000111011101),
      .k8(32'b00111110000100011000101001111010),
      .k9(32'b00111110000111000111011000100101)
  ) CON2D_94(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[31]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101101011110110010100001110),
      .k2(32'b00111101110000110001010100010101),
      .k3(32'b00111110000001010111111001000010),
      .k4(32'b10111100011011101110101010011100),
      .k5(32'b00111011101011110101000111110101),
      .k6(32'b00111101001011001100110101001110),
      .k7(32'b00111101110000100111011111111011),
      .k8(32'b00111101101110001110110010101001),
      .k9(32'b00111101111001000110010110111010)
  ) CON2D_95(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[31]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111110001001000011000001),
      .k2(32'b00111101111001000010110000111110),
      .k3(32'b00111110000010010101111011100000),
      .k4(32'b00111101111000110101101001001101),
      .k5(32'b00111101111000011010101100101011),
      .k6(32'b00111110000010000100111011100111),
      .k7(32'b00111110000111011010101111101110),
      .k8(32'b00111110000001000011100100100011),
      .k9(32'b00111110000011001101011000011000)
  ) CON2D_96(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[31]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op31(
      .o_CORE_IP1(o_CORE_IP1[31]), 
      .o_CORE_IP2(o_CORE_IP2[31]), 
      .o_CORE_IP3(o_CORE_IP3[31]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data31), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111000101000001000011111),
      .k2(32'b10111101100110001101010101001111),
      .k3(32'b00111100010110010100100010101000),
      .k4(32'b10111101101111010100010111000001),
      .k5(32'b10111101010000101000110001011111),
      .k6(32'b00111101011101000001101000110011),
      .k7(32'b10111101110100101001101001110001),
      .k8(32'b10111101100101001000010011110111),
      .k9(32'b00111100001100100110111111011011)
  ) CON2D_97(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[32]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111111010100100110110000),
      .k2(32'b10111101101000000110000101010110),
      .k3(32'b00111101000001101101111010111100),
      .k4(32'b10111101100000011111111000001000),
      .k5(32'b10111011111011100111000101001111),
      .k6(32'b00111101111111000101110110110100),
      .k7(32'b10111101110100000111011101110110),
      .k8(32'b10111101011110000010111010001001),
      .k9(32'b00111101001101111110011100010010)
  ) CON2D_98(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[32]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101110110101111011001111000),
      .k2(32'b10111101100100011111101010010010),
      .k3(32'b00111100100110110001110100100001),
      .k4(32'b10111101110110010010000000011010),
      .k5(32'b10111101011110110010101001000011),
      .k6(32'b00111101010001000100000101111110),
      .k7(32'b10111101110111000100110100111100),
      .k8(32'b10111101100111001010001101000110),
      .k9(32'b00111100000001011011011001101100)
  ) CON2D_99(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[32]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op32(
      .o_CORE_IP1(o_CORE_IP1[32]), 
      .o_CORE_IP2(o_CORE_IP2[32]), 
      .o_CORE_IP3(o_CORE_IP3[32]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data32), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111011101110110011011100100101),
      .k2(32'b10111110000111111101111001011001),
      .k3(32'b10111011101001001111001101000010),
      .k4(32'b00111110010001011100000110010010),
      .k5(32'b00111101001001010100000111010000),
      .k6(32'b00111110001111001010001001100011),
      .k7(32'b00111101111011110000101110111010),
      .k8(32'b10111100110010000011000111011101),
      .k9(32'b00111101111100111110111010111011)
  ) CON2D_100(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[33]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111100100101001110011001000000),
      .k2(32'b10111110010010100100010011010100),
      .k3(32'b10111101000110011000110011011111),
      .k4(32'b00111110100100010010100001101110),
      .k5(32'b00111101111011001000001011001100),
      .k6(32'b00111110100001111110000100100011),
      .k7(32'b00111110010100110000001001011111),
      .k8(32'b00111101010101001110011011100011),
      .k9(32'b00111110010010110100111001111000)
  ) CON2D_101(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[33]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111110011010011111111100),
      .k2(32'b10111110100111101101101000100111),
      .k3(32'b10111110000110001011000110011011),
      .k4(32'b10111100101100000011000101110100),
      .k5(32'b10111110010100000001001011111011),
      .k6(32'b10111101001011010110011011101110),
      .k7(32'b10111100000100110010111010001000),
      .k8(32'b10111110001100101001000010111010),
      .k9(32'b10111100100111110000111010110110)
  ) CON2D_102(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[33]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op33(
      .o_CORE_IP1(o_CORE_IP1[33]), 
      .o_CORE_IP2(o_CORE_IP2[33]), 
      .o_CORE_IP3(o_CORE_IP3[33]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data33), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110011110101010101111110011),
      .k2(32'b10111110100101000111101101010110),
      .k3(32'b10111110100010100100011100010001),
      .k4(32'b00111101110000111010101100010100),
      .k5(32'b00111110000000100100110011001011),
      .k6(32'b00111101111010101111001001011001),
      .k7(32'b00111101101111111000101100000100),
      .k8(32'b00111110001010110101001001100000),
      .k9(32'b00111110000110001111010000101111)
  ) CON2D_103(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[34]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100001100111010111000000),
      .k2(32'b10111110101001001111101001111000),
      .k3(32'b10111110100110111010001101110001),
      .k4(32'b00111110101111110111110010011110),
      .k5(32'b00111110110011011001110010001111),
      .k6(32'b00111110110000011001011111001010),
      .k7(32'b00111110101110101111111001010010),
      .k8(32'b00111110111000001110100011100110),
      .k9(32'b00111110110100001000010101101111)
  ) CON2D_104(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[34]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110101011000011111111111101),
      .k2(32'b10111110110110101101111100101101),
      .k3(32'b10111110110011000000111000101010),
      .k4(32'b10111101101100101101110110111001),
      .k5(32'b10111101110110101100110111000100),
      .k6(32'b10111101110101000000101110110010),
      .k7(32'b10111011010010100111100011011110),
      .k8(32'b00111100110110101101100111011010),
      .k9(32'b00111100101111110001111101110100)
  ) CON2D_105(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[34]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op34(
      .o_CORE_IP1(o_CORE_IP1[34]), 
      .o_CORE_IP2(o_CORE_IP2[34]), 
      .o_CORE_IP3(o_CORE_IP3[34]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data34), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100111000101000010100111),
      .k2(32'b10111110110111010101000100111100),
      .k3(32'b10111110110011100111010000001001),
      .k4(32'b10111110011101110011100100110001),
      .k5(32'b10111110101001011110001011010010),
      .k6(32'b10111110100110111110011011001000),
      .k7(32'b10111101110101100100001001010110),
      .k8(32'b10111110000100111111100110111101),
      .k9(32'b10111110000011010100100000100100)
  ) CON2D_106(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[35]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001010111000111001001110),
      .k2(32'b10111110010100111011001010101011),
      .k3(32'b10111110010001110100100011101001),
      .k4(32'b00111110000100011011010001001000),
      .k5(32'b00111110001001110011011100110110),
      .k6(32'b00111110000111100000100111101111),
      .k7(32'b00111101110001110101111000010010),
      .k8(32'b00111110000110000110100101110101),
      .k9(32'b00111110000001011001110111000000)
  ) CON2D_107(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[35]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101000010110010011001010010),
      .k2(32'b00111101100110110100000011001010),
      .k3(32'b00111101100010010101001001001010),
      .k4(32'b00111110101100000011010011110010),
      .k5(32'b00111110111000111001001110001110),
      .k6(32'b00111110110100011000001010100000),
      .k7(32'b00111110001111101001001100101111),
      .k8(32'b00111110100110110011011000011101),
      .k9(32'b00111110100010000000101100010111)
  ) CON2D_108(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[35]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op35(
      .o_CORE_IP1(o_CORE_IP1[35]), 
      .o_CORE_IP2(o_CORE_IP2[35]), 
      .o_CORE_IP3(o_CORE_IP3[35]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data35), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101011110011001101000011111),
      .k2(32'b00111101010011110110001100011001),
      .k3(32'b10111110001011111100001001110100),
      .k4(32'b00111101100101011110001010010110),
      .k5(32'b00111101001010101011110100111001),
      .k6(32'b10111110010011111111001111110001),
      .k7(32'b00111101011111010110110111010010),
      .k8(32'b00111101010010011100100010111101),
      .k9(32'b10111110001100100101000011011110)
  ) CON2D_109(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[36]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101100011011001101010110001),
      .k2(32'b00111101001001111000011010111010),
      .k3(32'b10111110010100001011111010001011),
      .k4(32'b00111101101101101001110001101100),
      .k5(32'b00111101000111110100111100111001),
      .k6(32'b10111110011010011111101000010011),
      .k7(32'b00111101100110100101011100010010),
      .k8(32'b00111101001110000101010111110100),
      .k9(32'b10111110010011001001001010001000)
  ) CON2D_110(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[36]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101011101100101111101011110),
      .k2(32'b00111101010101010000100100101110),
      .k3(32'b10111110001100010011100010000010),
      .k4(32'b00111101100101111110101010101010),
      .k5(32'b00111101001101011011100111011111),
      .k6(32'b10111110010011111001110101000100),
      .k7(32'b00111101100010000100011101010000),
      .k8(32'b00111101011000000011010100111011),
      .k9(32'b10111110001011100101111101101100)
  ) CON2D_111(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[36]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op36(
      .o_CORE_IP1(o_CORE_IP1[36]), 
      .o_CORE_IP2(o_CORE_IP2[36]), 
      .o_CORE_IP3(o_CORE_IP3[36]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data36), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110101010000000010011101011),
      .k2(32'b10111110110111001011000001001101),
      .k3(32'b10111110101111001110000000101000),
      .k4(32'b10111101110011000001010011111111),
      .k5(32'b10111101111101101011001001101111),
      .k6(32'b10111101101100110001110011111010),
      .k7(32'b00111101001101101001101010101010),
      .k8(32'b00111101100111000000010001101101),
      .k9(32'b00111101100110100101101000110110)
  ) CON2D_112(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[37]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100011110100100011000001),
      .k2(32'b10111110101100110011100000001101),
      .k3(32'b10111110100100010100001101101001),
      .k4(32'b00111110101010110001000101000100),
      .k5(32'b00111110101110010100111000110001),
      .k6(32'b00111110110000110000101111101111),
      .k7(32'b00111110111010110100100100010111),
      .k8(32'b00111111000010100001101010011110),
      .k9(32'b00111111000001001011100010010000)
  ) CON2D_113(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[37]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100101111001101010001010),
      .k2(32'b10111110101110010111011110110011),
      .k3(32'b10111110100110000010100011100101),
      .k4(32'b00111011100101001010010111010001),
      .k5(32'b00111100101111110100000010010000),
      .k6(32'b00111101010101111101010001010001),
      .k7(32'b00111110000010011101110011100000),
      .k8(32'b00111110010011101001000111100010),
      .k9(32'b00111110010010001100001010111100)
  ) CON2D_114(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[37]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op37(
      .o_CORE_IP1(o_CORE_IP1[37]), 
      .o_CORE_IP2(o_CORE_IP2[37]), 
      .o_CORE_IP3(o_CORE_IP3[37]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data37), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001011110100110111010010),
      .k2(32'b00111110100101101100000100010110),
      .k3(32'b00111110000001011111010001100000),
      .k4(32'b00111100100001101011101011100001),
      .k5(32'b00111101110011110100001111000011),
      .k6(32'b10111101100000000000110001000000),
      .k7(32'b10111101101101100000011001010010),
      .k8(32'b10111101000110001111101101110001),
      .k9(32'b10111110001011100011000100111000)
  ) CON2D_115(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[38]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110010111011110010111111101),
      .k2(32'b00111110101010001000111001001111),
      .k3(32'b00111110000111100100111001101111),
      .k4(32'b00111011100011001011101111000111),
      .k5(32'b00111101100101110010011101010101),
      .k6(32'b10111101110010011111000101000001),
      .k7(32'b10111110000001000111100110001001),
      .k8(32'b10111101110000111111110101010000),
      .k9(32'b10111110011100011000000101101011)
  ) CON2D_116(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[38]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101011001110110011000100110),
      .k2(32'b00111110000110100000011011101110),
      .k3(32'b10111010101011101000111011101111),
      .k4(32'b10111101101011000011000001110100),
      .k5(32'b10111100111111101110100110010001),
      .k6(32'b10111110001110111001000101010000),
      .k7(32'b10111110000010010010100100001100),
      .k8(32'b10111101111000111001100001000011),
      .k9(32'b10111110011100000010110010100001)
  ) CON2D_117(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[38]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op38(
      .o_CORE_IP1(o_CORE_IP1[38]), 
      .o_CORE_IP2(o_CORE_IP2[38]), 
      .o_CORE_IP3(o_CORE_IP3[38]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data38), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110100100011110001001100),
      .k2(32'b10111101111000010010011010001110),
      .k3(32'b10111101000100101111111110000001),
      .k4(32'b00111101111110000011100101000010),
      .k5(32'b10111101111010000010111100111011),
      .k6(32'b10111101001010111110100101001110),
      .k7(32'b00111101110100010110000001010110),
      .k8(32'b10111101110101010100011100100101),
      .k9(32'b10111101000001010111100101001110)
  ) CON2D_118(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[39]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001111000011101100101011),
      .k2(32'b10111110010010100101010000111100),
      .k3(32'b10111101111101011001000000110111),
      .k4(32'b00111100100110101000100000001010),
      .k5(32'b10111110011111101101010001011001),
      .k6(32'b10111110001100010110101111000101),
      .k7(32'b00111101010001110001001110110000),
      .k8(32'b10111110001111101110101000101000),
      .k9(32'b10111101111000110111000101110111)
  ) CON2D_119(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[39]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101101110011011010011101000),
      .k2(32'b10111110000000000110001111001011),
      .k3(32'b10111101001111100011010110111111),
      .k4(32'b00111101110011110001110111010101),
      .k5(32'b10111110000010111001101110011001),
      .k6(32'b10111101011101000110001110000001),
      .k7(32'b00111101101001001000101100101101),
      .k8(32'b10111110000000101111111011111111),
      .k9(32'b10111101010100011011111100101100)
  ) CON2D_120(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[39]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op39(
      .o_CORE_IP1(o_CORE_IP1[39]), 
      .o_CORE_IP2(o_CORE_IP2[39]), 
      .o_CORE_IP3(o_CORE_IP3[39]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data39), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111000101001010101111000),
      .k2(32'b00111101100001111010010111011110),
      .k3(32'b10111101110110011010000001101111),
      .k4(32'b10111100100101100101101111110100),
      .k5(32'b00111110010001110010100110000010),
      .k6(32'b10111010101000010111001011100111),
      .k7(32'b10111101001001111000011111101100),
      .k8(32'b00111110001100010111110011111000),
      .k9(32'b10111100011001010000011101101110)
  ) CON2D_121(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[40]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111001100100010010011101),
      .k2(32'b00111101100001101101110010000000),
      .k3(32'b10111101111010101000110100011111),
      .k4(32'b00111100110010000000001010101010),
      .k5(32'b00111110011101100000000000011100),
      .k6(32'b00111101000100011110110010101000),
      .k7(32'b10111100100001010101110111110110),
      .k8(32'b00111110010011011111111111101001),
      .k9(32'b00111011101011000010100100001010)
  ) CON2D_122(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[40]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000111110110110001000101),
      .k2(32'b10111011100000110110110000111010),
      .k3(32'b10111110001001111010011111110100),
      .k4(32'b10111101110101011111011010001011),
      .k5(32'b00111101101000001100011010001101),
      .k6(32'b10111101110100101001000110100010),
      .k7(32'b10111101110110101010010111111111),
      .k8(32'b00111101101000011010110110000100),
      .k9(32'b10111101110000100101111101010100)
  ) CON2D_123(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[40]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op40(
      .o_CORE_IP1(o_CORE_IP1[40]), 
      .o_CORE_IP2(o_CORE_IP2[40]), 
      .o_CORE_IP3(o_CORE_IP3[40]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data40), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101010010000011011001000),
      .k2(32'b00111110001110001001111110000011),
      .k3(32'b00111110100101010010111001110000),
      .k4(32'b10111011100100100110100010111111),
      .k5(32'b10111110011011010111000000010011),
      .k6(32'b10111101110001101111100110011111),
      .k7(32'b10111101111010011000100100111000),
      .k8(32'b10111110101110110011111010100000),
      .k9(32'b10111110011001000011111000100001)
  ) CON2D_124(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[41]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101101111100010100111000),
      .k2(32'b00111110010100000100100000011101),
      .k3(32'b00111110100111111001001110001010),
      .k4(32'b10111110001011010110011001101100),
      .k5(32'b10111110110100001001010100000001),
      .k6(32'b10111110100010100110000000100111),
      .k7(32'b10111110100100100101111001011000),
      .k8(32'b10111111000011010011111111001000),
      .k9(32'b10111110110011110010101101000010)
  ) CON2D_125(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[41]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110110010101101010110000101),
      .k2(32'b00111110100100010001110110000001),
      .k3(32'b00111110110000010011001001101001),
      .k4(32'b00111110010111101100100100000110),
      .k5(32'b00111101000111111001111000001101),
      .k6(32'b00111110000111000100011010000101),
      .k7(32'b00111101101100000100101010010110),
      .k8(32'b10111101111011011110011101111101),
      .k9(32'b00111011111110111010110100011000)
  ) CON2D_126(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[41]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op41(
      .o_CORE_IP1(o_CORE_IP1[41]), 
      .o_CORE_IP2(o_CORE_IP2[41]), 
      .o_CORE_IP3(o_CORE_IP3[41]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data41), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101011100000110110010010000),
      .k2(32'b10111101100100000110001000010110),
      .k3(32'b10111101100000010011111001001111),
      .k4(32'b10111110010000101100101000000101),
      .k5(32'b10111110011011000001100111110101),
      .k6(32'b10111110010111111101100010001100),
      .k7(32'b10111110010001000000011111100101),
      .k8(32'b10111110011111111011010110010110),
      .k9(32'b10111110011010110101000001101010)
  ) CON2D_127(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[42]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000011010000111011000000),
      .k2(32'b00111110001011010000011111110111),
      .k3(32'b00111110000110100000111000001010),
      .k4(32'b00111100101000110110001111000000),
      .k5(32'b00111100110011100111001010010001),
      .k6(32'b00111100010101011000110100011100),
      .k7(32'b10111110000001000011100101101101),
      .k8(32'b10111110000111000100110110110010),
      .k9(32'b10111110000110001101011001101101)
  ) CON2D_128(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[42]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011000101100000001000101),
      .k2(32'b00111110100100100001110010111000),
      .k3(32'b00111110100000010101010111010111),
      .k4(32'b00111110010001111100101110100101),
      .k5(32'b00111110011101100110111010111000),
      .k6(32'b00111110010110000011110000111010),
      .k7(32'b00111001111110001010000111101100),
      .k8(32'b00111100011111110110011111010000),
      .k9(32'b00111011110000101110100100111000)
  ) CON2D_129(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[42]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op42(
      .o_CORE_IP1(o_CORE_IP1[42]), 
      .o_CORE_IP2(o_CORE_IP2[42]), 
      .o_CORE_IP3(o_CORE_IP3[42]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data42), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001111010011100011011001),
      .k2(32'b00111110100111011000110100110011),
      .k3(32'b00111110100100101001110111000110),
      .k4(32'b10111101100001000111010100000100),
      .k5(32'b10111101000000100101100000001101),
      .k6(32'b10111100101110001101000000101111),
      .k7(32'b10111101111000011001101010110000),
      .k8(32'b10111110000100110011001110110001),
      .k9(32'b10111101111101001000100000000010)
  ) CON2D_130(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[43]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110001110110101101000110111),
      .k2(32'b00111110100110001100010000110011),
      .k3(32'b00111110100011100111010110010000),
      .k4(32'b10111110101010011101011111100000),
      .k5(32'b10111110101001010010011010101100),
      .k6(32'b10111110100111010011010011111100),
      .k7(32'b10111110110000101000110110001100),
      .k8(32'b10111110111000110010010011101111),
      .k9(32'b10111110110100101111001111010001)
  ) CON2D_131(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[43]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110010110100101100000001110),
      .k2(32'b00111110101011101011101101010010),
      .k3(32'b00111110100111011110100101111001),
      .k4(32'b10111100011010001011010100001101),
      .k5(32'b00111100110110000010100110001111),
      .k6(32'b00111100110010001100010000101101),
      .k7(32'b10111101101101110100000100110110),
      .k8(32'b10111101111011110010001010000000),
      .k9(32'b10111101110100101110101010101010)
  ) CON2D_132(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[43]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op43(
      .o_CORE_IP1(o_CORE_IP1[43]), 
      .o_CORE_IP2(o_CORE_IP2[43]), 
      .o_CORE_IP3(o_CORE_IP3[43]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data43), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100001011000010101111110100),
      .k2(32'b00111101110001100000100100010101),
      .k3(32'b10111101001011100100011101100101),
      .k4(32'b00111110001011110000111101011111),
      .k5(32'b00111110100011110010111101101101),
      .k6(32'b00111101111011110111000000111100),
      .k7(32'b00111101100011000110111010001100),
      .k8(32'b00111110001111000000100111100000),
      .k9(32'b00111101000100011001101000000010)
  ) CON2D_133(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[44]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101011000100000010010110100),
      .k2(32'b00111011100110010011110100001110),
      .k3(32'b10111110000001111101000001100010),
      .k4(32'b00111110000011100001010111101011),
      .k5(32'b00111110011000101100100110101100),
      .k6(32'b00111101011110110110011001111101),
      .k7(32'b00111101011010111010000101110100),
      .k8(32'b00111110000110001111101000101011),
      .k9(32'b00111010101110000111100100101001)
  ) CON2D_134(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[44]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001101000111111011011101),
      .k2(32'b10111110000110100000010101100011),
      .k3(32'b10111110100000110011110001111100),
      .k4(32'b10111110000010000111110001100110),
      .k5(32'b10111101101110110101100001101100),
      .k6(32'b10111110010111000000100000101110),
      .k7(32'b10111101111010101111000110001110),
      .k8(32'b10111101011100110101010010011100),
      .k9(32'b10111110001100100110000011111110)
  ) CON2D_135(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[44]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op44(
      .o_CORE_IP1(o_CORE_IP1[44]), 
      .o_CORE_IP2(o_CORE_IP2[44]), 
      .o_CORE_IP3(o_CORE_IP3[44]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data44), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110110100111101100101111),
      .k2(32'b00111101110010100110110010011111),
      .k3(32'b00111101110100111101111011011011),
      .k4(32'b10111110110000010001001001111001),
      .k5(32'b10111110111101100000111011101100),
      .k6(32'b10111110111000011111000011001100),
      .k7(32'b10111110101011100110111100111110),
      .k8(32'b10111110111110001101110000111010),
      .k9(32'b10111110111000000011101000011100)
  ) CON2D_136(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[45]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100100101000110100100101),
      .k2(32'b00111110101101100110010110000011),
      .k3(32'b00111110101010010011001010100011),
      .k4(32'b10111110011110111001110110110000),
      .k5(32'b10111110100001111010010010100001),
      .k6(32'b10111110100000000101100100101010),
      .k7(32'b10111110100101110101011101110010),
      .k8(32'b10111110101111000111000111011001),
      .k9(32'b10111110101011010011101101101100)
  ) CON2D_137(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[45]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110110110011010011111011111),
      .k2(32'b00111111000100110011101001100011),
      .k3(32'b00111111000000110101000000101101),
      .k4(32'b00111110100111010100010100001110),
      .k5(32'b00111110110010111000110101100100),
      .k6(32'b00111110101110100110110011101000),
      .k7(32'b00111110000001110110111000010110),
      .k8(32'b00111110001010110111010000100000),
      .k9(32'b00111110001000000011000011011110)
  ) CON2D_138(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[45]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op45(
      .o_CORE_IP1(o_CORE_IP1[45]), 
      .o_CORE_IP2(o_CORE_IP2[45]), 
      .o_CORE_IP3(o_CORE_IP3[45]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data45), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000001100000001010010110),
      .k2(32'b10111101100010011100010001000101),
      .k3(32'b10111100111010010101010110100011),
      .k4(32'b00111101010110110101000100000110),
      .k5(32'b00111110001111101111110111100110),
      .k6(32'b00111110011001101110110100111100),
      .k7(32'b10111100100011000101100000111000),
      .k8(32'b00111101111011010101010101010101),
      .k9(32'b00111110000100110011110111110101)
  ) CON2D_139(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[46]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001111110011100101011001),
      .k2(32'b10111110000010101000110000110101),
      .k3(32'b10111101100110111010101000001110),
      .k4(32'b00111101111100000010110010100110),
      .k5(32'b00111110011110011001110110000100),
      .k6(32'b00111110100110101010000000010110),
      .k7(32'b00111101001110001000101111010101),
      .k8(32'b00111110001100110111111001010010),
      .k9(32'b00111110011000010001100011011000)
  ) CON2D_140(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[46]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100000011100101111010010),
      .k2(32'b10111110100001000101110001011110),
      .k3(32'b10111110010011101000001001001100),
      .k4(32'b10111110001110000100001100000101),
      .k5(32'b10111101111111111111100111110101),
      .k6(32'b10111101011101100100101110110011),
      .k7(32'b10111110000101001100111111101111),
      .k8(32'b10111101101001010010010111110010),
      .k9(32'b10111101000000011001110000000010)
  ) CON2D_141(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[46]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op46(
      .o_CORE_IP1(o_CORE_IP1[46]), 
      .o_CORE_IP2(o_CORE_IP2[46]), 
      .o_CORE_IP3(o_CORE_IP3[46]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data46), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110101110011100011000011000),
      .k2(32'b10111110111101111101011001010101),
      .k3(32'b10111110111001110001110111000110),
      .k4(32'b10111110001111011011000101111001),
      .k5(32'b10111110011100010110001010010110),
      .k6(32'b10111110011000101111000101010100),
      .k7(32'b00111101111010111011110110101101),
      .k8(32'b00111110000111011010000001101011),
      .k9(32'b00111110000100100111100010111100)
  ) CON2D_142(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[47]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110110000111101010011000011),
      .k2(32'b10111110111011100110001010001010),
      .k3(32'b10111110111000110001110010111111),
      .k4(32'b10111100000001010111001101110100),
      .k5(32'b10111011101000100001000010101010),
      .k6(32'b10111100001101110011110101100011),
      .k7(32'b00111110101100000110101011000001),
      .k8(32'b00111110110111110011001011110111),
      .k9(32'b00111110110011000010101110010101)
  ) CON2D_143(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[47]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101100101100111110011101000),
      .k2(32'b10111101101110011110011111010100),
      .k3(32'b10111101101100101000100110010001),
      .k4(32'b00111110010101110100110111011011),
      .k5(32'b00111110100010100010011000111000),
      .k6(32'b00111110011110011000111110100100),
      .k7(32'b00111110101001101110000010101110),
      .k8(32'b00111110111010001110001100100110),
      .k9(32'b00111110110100000110110000010110)
  ) CON2D_144(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[47]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op47(
      .o_CORE_IP1(o_CORE_IP1[47]), 
      .o_CORE_IP2(o_CORE_IP2[47]), 
      .o_CORE_IP3(o_CORE_IP3[47]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data47), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101100000111110100001100001),
      .k2(32'b00111110001010111001011001000110),
      .k3(32'b00111110010010001110010011011101),
      .k4(32'b00111110001001011101110110110111),
      .k5(32'b00111110100111011011101000001100),
      .k6(32'b00111110101011100110010110001000),
      .k7(32'b00111101100111110110101101010001),
      .k8(32'b00111110011100000100101110010000),
      .k9(32'b00111110100000110001000110001011)
  ) CON2D_145(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[48]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101110101000011101011011001),
      .k2(32'b10111101101111010110010011010111),
      .k3(32'b10111101000101111000101011011100),
      .k4(32'b10111100111101010011001000001111),
      .k5(32'b00111100101011110000110001001111),
      .k6(32'b00111101101011000000010011110110),
      .k7(32'b00111101011001110001100101101010),
      .k8(32'b00111110000010111110110010110010),
      .k9(32'b00111110001110001010100101011000)
  ) CON2D_146(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[48]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100001011110100101011000),
      .k2(32'b10111110101101110100011111001110),
      .k3(32'b10111110100110100111110000011010),
      .k4(32'b10111110101010010001111100101110),
      .k5(32'b10111110110011000001010001001000),
      .k6(32'b10111110101010010101000001000101),
      .k7(32'b10111101111000011101100001000011),
      .k8(32'b10111110000010100000000111000010),
      .k9(32'b10111101101100111011101111010010)
  ) CON2D_147(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[48]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op48(
      .o_CORE_IP1(o_CORE_IP1[48]), 
      .o_CORE_IP2(o_CORE_IP2[48]), 
      .o_CORE_IP3(o_CORE_IP3[48]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data48), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101101111110011001101100001),
      .k2(32'b10111101011000100100100000101011),
      .k3(32'b10111101101101111110010101111000),
      .k4(32'b10111110001001011000001101111100),
      .k5(32'b10111110101110101100110001000110),
      .k6(32'b10111110110011101101100001010000),
      .k7(32'b10111110000011000011101000110110),
      .k8(32'b10111110101010011001100101011100),
      .k9(32'b10111110101100110101100111011001)
  ) CON2D_148(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[49]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110100001100000111101100100),
      .k2(32'b00111110000010100000000011100011),
      .k3(32'b00111101011100000101000100101110),
      .k4(32'b00111100101111010100101000100111),
      .k5(32'b10111110000111101111100000111111),
      .k6(32'b10111110011100011100111101101111),
      .k7(32'b00111100011100101011101010011100),
      .k8(32'b10111110001000110111011001100011),
      .k9(32'b10111110010111100011000101010011)
  ) CON2D_149(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[49]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110110010110010000010001100),
      .k2(32'b00111110101010101001111110100101),
      .k3(32'b00111110100000011010011111111111),
      .k4(32'b00111110101011010010010100001111),
      .k5(32'b00111110011011110001111011011100),
      .k6(32'b00111110000100101000000010001101),
      .k7(32'b00111110011010101001110111010010),
      .k8(32'b00111101111111111011110111111111),
      .k9(32'b00111101011110010101100010100000)
  ) CON2D_150(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[49]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op49(
      .o_CORE_IP1(o_CORE_IP1[49]), 
      .o_CORE_IP2(o_CORE_IP2[49]), 
      .o_CORE_IP3(o_CORE_IP3[49]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data49), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111011100000111001101001000100),
      .k2(32'b00111110000000001010110100011011),
      .k3(32'b10111110000110101011110011001111),
      .k4(32'b00111100101010010001001000010011),
      .k5(32'b00111110000011100100011010111000),
      .k6(32'b10111110001000100001100100010000),
      .k7(32'b00111011101000110011000001110011),
      .k8(32'b00111101111111110100110111100011),
      .k9(32'b10111110000111100000001001000101)
  ) CON2D_151(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[50]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100001010001110111011101101),
      .k2(32'b00111110000010011100000011000010),
      .k3(32'b10111110001001011111110011101001),
      .k4(32'b00111101001011010100111000000101),
      .k5(32'b00111110001001101000100110010001),
      .k6(32'b10111110000111101001001110110010),
      .k7(32'b00111100100001001010111010001010),
      .k8(32'b00111110000011000000011011111011),
      .k9(32'b10111110001001010100000100000011)
  ) CON2D_152(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[50]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111011100001101110010111000111),
      .k2(32'b00111110000001111100111101010101),
      .k3(32'b10111110000101100100101011101100),
      .k4(32'b00111100101100001011101011101001),
      .k5(32'b00111110000101001111111010100111),
      .k6(32'b10111110000111011111111000011011),
      .k7(32'b00111100001010111110000111110010),
      .k8(32'b00111110000010001110111111011000),
      .k9(32'b10111110000101101010111101001100)
  ) CON2D_153(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[50]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op50(
      .o_CORE_IP1(o_CORE_IP1[50]), 
      .o_CORE_IP2(o_CORE_IP2[50]), 
      .o_CORE_IP3(o_CORE_IP3[50]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data50), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110110000011001110010011111),
      .k2(32'b00111111000000000001101001000111),
      .k3(32'b00111110111011010110101000100110),
      .k4(32'b00111110101010100111100101001010),
      .k5(32'b00111110110110011000110111000110),
      .k6(32'b00111110110010111101110001010111),
      .k7(32'b00111110100010101011100011110000),
      .k8(32'b00111110101101111001001100111111),
      .k9(32'b00111110101001111100011001110001)
  ) CON2D_154(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[51]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110000110011000111010100111),
      .k2(32'b00111110001000011011100100010000),
      .k3(32'b00111110001010100000000101100101),
      .k4(32'b10111110011000011110010111111011),
      .k5(32'b10111110100010000101001001100011),
      .k6(32'b10111110011101100110110010101101),
      .k7(32'b10111100001111111111110101100111),
      .k8(32'b10111101001110000010111101011000),
      .k9(32'b10111101000000110011011000010011)
  ) CON2D_155(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[51]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101110010111000100100010101),
      .k2(32'b10111110010000001111101000011000),
      .k3(32'b10111110000101100100001111010010),
      .k4(32'b10111111000001001100100110110001),
      .k5(32'b10111111001010111110000011100000),
      .k6(32'b10111111000111001011101101001111),
      .k7(32'b10111110011001000111001111100000),
      .k8(32'b10111110101100110111111001000101),
      .k9(32'b10111110100111100001110000101001)
  ) CON2D_156(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[51]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op51(
      .o_CORE_IP1(o_CORE_IP1[51]), 
      .o_CORE_IP2(o_CORE_IP2[51]), 
      .o_CORE_IP3(o_CORE_IP3[51]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data51), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101010101111100111101101010),
      .k2(32'b10111101100110000110110101010011),
      .k3(32'b00111110000000100000101011011100),
      .k4(32'b10111101101001000011111111000111),
      .k5(32'b10111110011011101010111101111011),
      .k6(32'b10111010101000001110100001101000),
      .k7(32'b00111011000000001110000010000010),
      .k8(32'b10111110001000001010100101000000),
      .k9(32'b00111101000100101000010110001001)
  ) CON2D_157(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[52]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100110100000001111100001110),
      .k2(32'b10111101100111101101111000101100),
      .k3(32'b00111110001011001111110101101010),
      .k4(32'b10111110000110100001000111101010),
      .k5(32'b10111110100011100101100001101000),
      .k6(32'b00111010001101011000000110011101),
      .k7(32'b10111101010000100010111110000100),
      .k8(32'b10111110001110110001010011000110),
      .k9(32'b00111101010111011010010011100001)
  ) CON2D_158(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[52]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101101101001010001111101111),
      .k2(32'b00111100011110010000111001000100),
      .k3(32'b00111110011100111011111110010101),
      .k4(32'b00111101001010011110111010100111),
      .k5(32'b10111101001111000110000101011000),
      .k6(32'b00111110010100100000001000010000),
      .k7(32'b00111101011001110011011101110000),
      .k8(32'b10111101001011100101100101001110),
      .k9(32'b00111110001011011011101000110111)
  ) CON2D_159(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[52]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op52(
      .o_CORE_IP1(o_CORE_IP1[52]), 
      .o_CORE_IP2(o_CORE_IP2[52]), 
      .o_CORE_IP3(o_CORE_IP3[52]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data52), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100010101010010011100111),
      .k2(32'b10111110101011010110110011111111),
      .k3(32'b10111110100011000100011001101010),
      .k4(32'b10111110001000101011000011011111),
      .k5(32'b10111110000100101111011100001010),
      .k6(32'b10111101100100011101011010111000),
      .k7(32'b10111011101100010100000001001010),
      .k8(32'b00111101100100110110011010011101),
      .k9(32'b00111101111110110100011111110010)
  ) CON2D_160(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[53]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110101000010010101100101110),
      .k2(32'b10111110101010001011001011011101),
      .k3(32'b10111110100001101101000010011000),
      .k4(32'b10111110000010110000101000000010),
      .k5(32'b10111101011010010001110010110110),
      .k6(32'b00111100010100110001000110010101),
      .k7(32'b00111101000000010110001011000011),
      .k8(32'b00111110001011100010100100000100),
      .k9(32'b00111110010111101111010101111111)
  ) CON2D_161(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[53]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111011101110000110110000101100),
      .k2(32'b00111101000111110000110100100111),
      .k3(32'b00111101100011010011010101111000),
      .k4(32'b00111110000100010001000110011011),
      .k5(32'b00111110100010111001101010100101),
      .k6(32'b00111110100110111001000101010110),
      .k7(32'b00111101111001000101000111100001),
      .k8(32'b00111110100100001101101101011100),
      .k9(32'b00111110100110011001000100111011)
  ) CON2D_162(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[53]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op53(
      .o_CORE_IP1(o_CORE_IP1[53]), 
      .o_CORE_IP2(o_CORE_IP2[53]), 
      .o_CORE_IP3(o_CORE_IP3[53]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data53), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111000101000011000100011),
      .k2(32'b10111100110101100000111011001111),
      .k3(32'b00111101001110010000100100100010),
      .k4(32'b00111110100000011100100010101000),
      .k5(32'b00111110000010100011111001101000),
      .k6(32'b00111110010010001010011000011010),
      .k7(32'b00111110101001110101101000010001),
      .k8(32'b00111110011111010111011110011100),
      .k9(32'b00111110100110011110101110111101)
  ) CON2D_163(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[54]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000100111010001001000011),
      .k2(32'b10111110101010100110010010011000),
      .k3(32'b10111110011110110110001110110010),
      .k4(32'b10111101000011000100110000110111),
      .k5(32'b10111110010100000010101000101111),
      .k6(32'b10111101111111001011110111010010),
      .k7(32'b00111110011100010110101110010100),
      .k8(32'b00111101111100001010001101100100),
      .k9(32'b00111110001110111010011101001010)
  ) CON2D_164(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[54]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001011001000000110110000),
      .k2(32'b10111110101111000100011100100010),
      .k3(32'b10111110100010111101111110001101),
      .k4(32'b10111101101001100101110011011011),
      .k5(32'b10111110100001111001110001101110),
      .k6(32'b10111110001100110001101001011100),
      .k7(32'b00111110000111011101001011011010),
      .k8(32'b00111100101101010010000100111001),
      .k9(32'b00111101110011001011110011101001)
  ) CON2D_165(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[54]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op54(
      .o_CORE_IP1(o_CORE_IP1[54]), 
      .o_CORE_IP2(o_CORE_IP2[54]), 
      .o_CORE_IP3(o_CORE_IP3[54]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data54), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101111100100001000001011011),
      .k2(32'b10111101100101101001010110000110),
      .k3(32'b10111110011101000011011110011001),
      .k4(32'b10111101110010100100111100110110),
      .k5(32'b10111101001100010101001101110000),
      .k6(32'b10111110011010010011100110010101),
      .k7(32'b10111101000011010110001000010010),
      .k8(32'b00111101001010110010010110111011),
      .k9(32'b10111110000010001111110111001110)
  ) CON2D_166(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[55]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101010000010011111011100110),
      .k2(32'b00111100101010101010111011011100),
      .k3(32'b10111110001100110010110011011000),
      .k4(32'b00111100011000111100001000110011),
      .k5(32'b00111101110000110010011101000011),
      .k6(32'b10111101111110101100111111000010),
      .k7(32'b00111101010100001100101101000101),
      .k8(32'b00111110000110011100110111011010),
      .k9(32'b10111101011010101111111111011101)
  ) CON2D_167(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[55]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101011001011010111100100111),
      .k2(32'b00111110000111001101001111110001),
      .k3(32'b10111101001011000110000010110100),
      .k4(32'b00111110000100101010000100111101),
      .k5(32'b00111110100000011101011001001001),
      .k6(32'b00111101000011110110001000010111),
      .k7(32'b00111101111111000011000111010101),
      .k8(32'b00111110011111000110001010011110),
      .k9(32'b00111101001001010001000101110011)
  ) CON2D_168(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[55]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op55(
      .o_CORE_IP1(o_CORE_IP1[55]), 
      .o_CORE_IP2(o_CORE_IP2[55]), 
      .o_CORE_IP3(o_CORE_IP3[55]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data55), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101001100000001010110011001),
      .k2(32'b10111101111011000011010110111011),
      .k3(32'b00111100000101010111100011011111),
      .k4(32'b10111110000000100000000100000001),
      .k5(32'b10111110100111100011111110001000),
      .k6(32'b10111110001010001110100101101010),
      .k7(32'b10111100100000010100110001101010),
      .k8(32'b10111110001110110111001000000000),
      .k9(32'b10111101010101110101110001101010)
  ) CON2D_169(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[56]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101110010011100111110011100),
      .k2(32'b10111101001001011011111111101010),
      .k3(32'b00111101101100101001101101010000),
      .k4(32'b10111101110101000100011000010001),
      .k5(32'b10111110100001110101011001101101),
      .k6(32'b10111101111011001001001100111011),
      .k7(32'b00111011100010110000011010100111),
      .k8(32'b10111110000101000011010011010111),
      .k9(32'b10111100000011100010000001100100)
  ) CON2D_170(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[56]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110011010101110101010011000),
      .k2(32'b00111110000001001100100000110011),
      .k3(32'b00111110011011100011110100100110),
      .k4(32'b00111110001111011110011111110101),
      .k5(32'b00111101100101000001001110000111),
      .k6(32'b00111110010001000101100111100110),
      .k7(32'b00111110001000101100000011100000),
      .k8(32'b00111101010100101000010111110000),
      .k9(32'b00111110001001101110000010110001)
  ) CON2D_171(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[56]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op56(
      .o_CORE_IP1(o_CORE_IP1[56]), 
      .o_CORE_IP2(o_CORE_IP2[56]), 
      .o_CORE_IP3(o_CORE_IP3[56]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data56), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111110101101001101101101100001),
      .k2(32'b00111110001011101011100111101010),
      .k3(32'b00111110100110010110111101101000),
      .k4(32'b00111110100110010000010100010010),
      .k5(32'b00111101101111011101110101111111),
      .k6(32'b00111110011010111111110000010010),
      .k7(32'b00111110101001100110101000110111),
      .k8(32'b00111110000101100100100001010111),
      .k9(32'b00111110100011010010110100101111)
  ) CON2D_172(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[57]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111100001100010111110001),
      .k2(32'b10111110000010000101110011011000),
      .k3(32'b00111100110000111100101010011000),
      .k4(32'b10111110000000111100010101011111),
      .k5(32'b10111110110100110000101001111111),
      .k6(32'b10111110011101111100011011111011),
      .k7(32'b00111110000001001010000100100011),
      .k8(32'b10111101111010001101111000110110),
      .k9(32'b00111101001010000111010101100001)
  ) CON2D_173(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[57]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100101010000101100000001011),
      .k2(32'b10111110011111110110111110000000),
      .k3(32'b10111101101010110000100010000111),
      .k4(32'b10111110001111110010000111010111),
      .k5(32'b10111110111110101100001001001111),
      .k6(32'b10111110100111110101000111111110),
      .k7(32'b00111101010111001010000001000010),
      .k8(32'b10111110010100101001001010110011),
      .k9(32'b10111101001100010101111001011011)
  ) CON2D_174(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[57]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op57(
      .o_CORE_IP1(o_CORE_IP1[57]), 
      .o_CORE_IP2(o_CORE_IP2[57]), 
      .o_CORE_IP3(o_CORE_IP3[57]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data57), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100100011100000111001010),
      .k2(32'b10111110101111000010110001110000),
      .k3(32'b10111110101000111101010110011000),
      .k4(32'b10111110100100100110101000001100),
      .k5(32'b10111110101110010110101000111101),
      .k6(32'b10111110101000100101000100001010),
      .k7(32'b10111110100110100001101111111110),
      .k8(32'b10111110110010001010011100000000),
      .k9(32'b10111110101101010010111000110001)
  ) CON2D_175(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[58]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101001101011110000110111011),
      .k2(32'b10111101001001111010101010111011),
      .k3(32'b10111100111011010101110000110100),
      .k4(32'b00111110100011000000101100101101),
      .k5(32'b00111110100110000101110000010100),
      .k6(32'b00111110100101100001101100101111),
      .k7(32'b10111100101111111000000011001000),
      .k8(32'b10111100111000001010100111010101),
      .k9(32'b10111100110000111001100111001100)
  ) CON2D_176(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[58]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111101111001010011000101011110),
      .k2(32'b00111110001100011100000110000110),
      .k3(32'b00111110000110100111100100011011),
      .k4(32'b00111110111000111001110100100001),
      .k5(32'b00111111000001111000111111110100),
      .k6(32'b00111110111110001111010101110101),
      .k7(32'b00111101111100010000000011110011),
      .k8(32'b00111110001011110010011011010101),
      .k9(32'b00111110000100101100011111000001)
  ) CON2D_177(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[58]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op58(
      .o_CORE_IP1(o_CORE_IP1[58]), 
      .o_CORE_IP2(o_CORE_IP2[58]), 
      .o_CORE_IP3(o_CORE_IP3[58]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data58), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110010011111100001001101011),
      .k2(32'b00111110000010001001100011100001),
      .k3(32'b00111101101100101011010100111101),
      .k4(32'b10111110011111001100111110000101),
      .k5(32'b00111110001001000000010110000000),
      .k6(32'b00111110000110010111010110011101),
      .k7(32'b10111110010110110001000010001000),
      .k8(32'b00111110000100010110110000111110),
      .k9(32'b00111101111001011011110011101000)
  ) CON2D_178(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[59]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110011110101010111011001110),
      .k2(32'b00111110000100101011111000101110),
      .k3(32'b00111110000000000001101111101101),
      .k4(32'b10111110100100101101000000000011),
      .k5(32'b00111110001101000011110110011000),
      .k6(32'b00111110010001111001011010110111),
      .k7(32'b10111110100000101111010011000110),
      .k8(32'b00111110000111011011110001101100),
      .k9(32'b00111110000111010111011011001110)
  ) CON2D_179(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[59]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110010001100000011111011011),
      .k2(32'b00111110000010010000111011001011),
      .k3(32'b00111101101011110010011100100010),
      .k4(32'b10111110011100011100010101010101),
      .k5(32'b00111110001001011110010000111001),
      .k6(32'b00111110000110010111001010001110),
      .k7(32'b10111110010100110000001110101011),
      .k8(32'b00111110000100010011111000110101),
      .k9(32'b00111101111000011101101101011011)
  ) CON2D_180(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[59]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op59(
      .o_CORE_IP1(o_CORE_IP1[59]), 
      .o_CORE_IP2(o_CORE_IP2[59]), 
      .o_CORE_IP3(o_CORE_IP3[59]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data59), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100100011110010000101110),
      .k2(32'b10111110101110111101100110111000),
      .k3(32'b10111110101011010100110110111101),
      .k4(32'b10111110011010100111111101110010),
      .k5(32'b10111110100011010100100100010111),
      .k6(32'b10111110100001010100110001111011),
      .k7(32'b10111110001001100101100001010011),
      .k8(32'b10111110001110100110111001111111),
      .k9(32'b10111110001011110101000111010000)
  ) CON2D_181(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[60]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110001110010110000100011110),
      .k2(32'b10111110010100000001010111110011),
      .k3(32'b10111110010011101011111010111001),
      .k4(32'b00111110000100011000111110100010),
      .k5(32'b00111110001011001001011010101111),
      .k6(32'b00111110000100111001111111001110),
      .k7(32'b00111101101000110010011110000011),
      .k8(32'b00111110000000000011100001011001),
      .k9(32'b00111101110011110000001011000100)
  ) CON2D_182(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[60]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111100101000001101001000100100),
      .k2(32'b00111101010101010101010110100000),
      .k3(32'b00111101000010001010100011001011),
      .k4(32'b00111110101111010001100010110000),
      .k5(32'b00111110111001011111011101001010),
      .k6(32'b00111110110011001000111001001110),
      .k7(32'b00111110010101101000110111011011),
      .k8(32'b00111110100110010111100010001011),
      .k9(32'b00111110100000111000100000001011)
  ) CON2D_183(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[60]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op60(
      .o_CORE_IP1(o_CORE_IP1[60]), 
      .o_CORE_IP2(o_CORE_IP2[60]), 
      .o_CORE_IP3(o_CORE_IP3[60]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data60), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000001110110101001010110),
      .k2(32'b10111101101011011011011001100110),
      .k3(32'b10111110000000100010111111010011),
      .k4(32'b10111101111010100001111010010111),
      .k5(32'b10111101100011100000001100100001),
      .k6(32'b10111101110010100110110000000101),
      .k7(32'b10111110000100001101100000011100),
      .k8(32'b10111101110101110001001101001001),
      .k9(32'b10111110000110010101011000101000)
  ) CON2D_184(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[61]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000101111100001110011100),
      .k2(32'b10111101110010100111000111001111),
      .k3(32'b10111101111110101001100000101110),
      .k4(32'b10111101010101010000011101011001),
      .k5(32'b10111011011110000101111001001001),
      .k6(32'b10111100011001100111000011001001),
      .k7(32'b10111101111110110101100100101101),
      .k8(32'b10111101101010011100100010111011),
      .k9(32'b10111101111000001101010001100010)
  ) CON2D_185(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[61]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110000011111000010110101101),
      .k2(32'b10111101110000010010011011100000),
      .k3(32'b10111110000001001000001010100001),
      .k4(32'b10111110000101010111001010111010),
      .k5(32'b10111101110100111111100100010011),
      .k6(32'b10111110000000001011010010000100),
      .k7(32'b10111110000111001100010000111010),
      .k8(32'b10111101111100100100101001110010),
      .k9(32'b10111110001000001001101010011101)
  ) CON2D_186(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[61]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op61(
      .o_CORE_IP1(o_CORE_IP1[61]), 
      .o_CORE_IP2(o_CORE_IP2[61]), 
      .o_CORE_IP3(o_CORE_IP3[61]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data61), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101010110101000001011101111),
      .k2(32'b10111101010100010111011100001010),
      .k3(32'b10111101010011100000011001111111),
      .k4(32'b00111110101110110010001000011001),
      .k5(32'b00111110110111111100110111001000),
      .k6(32'b00111110110011101110000011000011),
      .k7(32'b00111110011101101110001011010011),
      .k8(32'b00111110101011011101100110000110),
      .k9(32'b00111110100111010001010100100100)
  ) CON2D_187(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[62]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110011100001111001010101000),
      .k2(32'b10111110100101111010011011111000),
      .k3(32'b10111110100011011000101011101000),
      .k4(32'b00111110100000111010100100001001),
      .k5(32'b00111110100010011111000001101101),
      .k6(32'b00111110100001001100001100010100),
      .k7(32'b00111110011110101000111101011001),
      .k8(32'b00111110100101110100011101010101),
      .k9(32'b00111110100011101111001111001011)
  ) CON2D_188(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[62]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110110000010101110110001011),
      .k2(32'b10111111000000010111001100011010),
      .k3(32'b10111110111011001010101100111000),
      .k4(32'b10111110100010110010110001110101),
      .k5(32'b10111110101100010000101110110010),
      .k6(32'b10111110101000001100100000001111),
      .k7(32'b10111110000011110100011001111101),
      .k8(32'b10111110001010110001000101000010),
      .k9(32'b10111110000100100100110110100100)
  ) CON2D_189(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[62]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op62(
      .o_CORE_IP1(o_CORE_IP1[62]), 
      .o_CORE_IP2(o_CORE_IP2[62]), 
      .o_CORE_IP3(o_CORE_IP3[62]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data62), 
      .valid_out()
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b00111011111110000100101110110100),
      .k2(32'b00111101000110011001001110101011),
      .k3(32'b00111101000011101110111110110100),
      .k4(32'b00111110101011100000110001111100),
      .k5(32'b00111110110100111000101100110101),
      .k6(32'b00111110110010001111110111001000),
      .k7(32'b00111101001110101001110101011001),
      .k8(32'b00111101110010100000001001101101),
      .k9(32'b00111101101101001100011011111110)
  ) CON2D_190(
      .i_data(o_fifo_in[31:0]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP1[63]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111101100000010001100011011010),
      .k2(32'b10111101100100000100000010011001),
      .k3(32'b10111101001000000001000111111100),
      .k4(32'b00111110101111100100110100110001),
      .k5(32'b00111110110100011010101011000010),
      .k6(32'b00111110110110001111011110101000),
      .k7(32'b00111101010110100100100000001100),
      .k8(32'b00111101100110000111011110101011),
      .k9(32'b00111101110000011101100100101111)
  ) CON2D_191(
      .i_data(o_fifo_in[63:32]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP2[63]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Con2D #(
      .DATA_WIDTH(DATA_WIDTH),
      .WIDTH(WIDTH+2),
      .k1(32'b10111110100110011101110001101110),
      .k2(32'b10111110110001000111001110010101),
      .k3(32'b10111110101001011110000101100110),
      .k4(32'b10111110011101010111100010101111),
      .k5(32'b10111110100101011100000011000010),
      .k6(32'b10111110011011100110110110001100),
      .k7(32'b10111110100001111011011111110001),
      .k8(32'b10111110101001001111110011100110),
      .k9(32'b10111110100010100001010101101010)
  ) CON2D_192(
      .i_data(o_fifo_in[95:64]),
      .valid_in(~empty_FIFO_IN),
      .clk(clk),
      .rst(rst),
      .fifo_busy(1'b0),
      .o_data(o_CORE_IP3[63]),
      .valid_out(),
      .rd_req(rd_req_FIFO_IN)
  );
  Op1_con3d#(
      .DATA_WIDTH(DATA_WIDTH),
      .bias(32'b00111111001110111111101011111010)
  )   op63(
      .o_CORE_IP1(o_CORE_IP1[63]), 
      .o_CORE_IP2(o_CORE_IP2[63]), 
      .o_CORE_IP3(o_CORE_IP3[63]), 
      .valid_in_adder(valid_in_adder), 
      .clk(clk), 
      .rst(rst), 
      .o_data(o_data63), 
      .valid_out()
  );
endmodule
