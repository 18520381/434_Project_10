module layer14_1#(
  parameter DATA_WIDTH = 32
  )(
  input  [DATA_WIDTH*32-1:0] i_data,
  input         clk, rst, valid_in,
  output [DATA_WIDTH*16-1:0] o_data ,
  output valid_out
  );
  
  wire [6:0] valid_pipeline_FC;

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110100101101111011010101101),
      .k2(32'b00111110100100110110011110001111),
      .k3(32'b00111110000011010000001111101100),
      .k4(32'b00111110011110110000010110011010),
      .k5(32'b00111110001011000010111100111110),
      .k6(32'b00111100101110100000010110000000),
      .k7(32'b00111101111100000110100100010100),
      .k8(32'b10111110101100001000011101110011),
      .k9(32'b10111110101010001001101010111010),
      .k10(32'b10111110100111011100010101101011),
      .k11(32'b00111110100000001011000000110101),
      .k12(32'b10111101100110011011010000101000),
      .k13(32'b10111101010110010001010110010000),
      .k14(32'b00111101010000100001011110011000),
      .k15(32'b00111100110000011011001011110000),
      .k16(32'b00111101100001110011101000001100),
      .k17(32'b10111101101010100111100011101000),
      .k18(32'b10111110001100101011101100110011),
      .k19(32'b00111100100101100110110111000000),
      .k20(32'b10111101110100101111000001111000),
      .k21(32'b10111110011001111010100110010011),
      .k22(32'b10111101110111110110000110001010),
      .k23(32'b00111110010111010000111110011110),
      .k24(32'b00111010000010111110011000000000),
      .k25(32'b10111101001110100001111001110000),
      .k26(32'b00111101100011100100110011110100),
      .k27(32'b10111101000001101001010011010000),
      .k28(32'b00111101010011110110001100011000),
      .k29(32'b10111110011111011000111110110010),
      .k30(32'b10111101110000001000110100110100),
      .k31(32'b10111110100111010101010111100101),
      .k32(32'b10111110100111010100011001111100),
      .bias(32'b00000000000000000000000000000000)
  ) FC1 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*1-1:DATA_WIDTH*0])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111101011001110101101001100001),
      .k2(32'b00111100111100110000111100111001),
      .k3(32'b10111110101010100011111011100010),
      .k4(32'b10111101101010110111110011010100),
      .k5(32'b10111110100010100011011110101100),
      .k6(32'b00111110100100111000100100101110),
      .k7(32'b00111110000001111010101111111101),
      .k8(32'b00111110010100111110101100111100),
      .k9(32'b00111110000011111000101100000010),
      .k10(32'b10111110001010010100100010100101),
      .k11(32'b10111110001010000011100001111011),
      .k12(32'b10111110011110011000111100000100),
      .k13(32'b10111110100101001011001111011001),
      .k14(32'b00111110100110000011100011000111),
      .k15(32'b10111110000110011010000110001110),
      .k16(32'b10111100100100010111010010101111),
      .k17(32'b00111100101011001011110101000110),
      .k18(32'b00111110000000110111000110101100),
      .k19(32'b10111110100101100101101000010011),
      .k20(32'b00111110001110010100010010010110),
      .k21(32'b00111100110100101001101011101101),
      .k22(32'b10111110101001111100111011101110),
      .k23(32'b00111110011011111110111000111100),
      .k24(32'b10111110100111010111101011011110),
      .k25(32'b10111110000110110010111100010110),
      .k26(32'b00111101101001100100111000001011),
      .k27(32'b10111110101011110111010101011111),
      .k28(32'b00111110100000001011001111010001),
      .k29(32'b10111101100101111110001110011001),
      .k30(32'b10111101111000000110110001110110),
      .k31(32'b00111110101011001101101111001000),
      .k32(32'b10111101100110111000000010100111),
      .bias(32'b00111011110101000010001111001110)
  ) FC2 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*2-1:DATA_WIDTH*1])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110101010001010100010000000),
      .k2(32'b10111101100000101001011100010001),
      .k3(32'b00111110100101100011010010111100),
      .k4(32'b00111110010011010100111011100011),
      .k5(32'b10111101100011110010001011101001),
      .k6(32'b00111110010101111101001110011000),
      .k7(32'b00111110011100110010110001101110),
      .k8(32'b00111110011110111110110001100100),
      .k9(32'b10111110101001110101100000100100),
      .k10(32'b00111110001010010101001011011001),
      .k11(32'b10111110000101001011100111000100),
      .k12(32'b10111110011110011010010010100110),
      .k13(32'b00111110000110111010110010001111),
      .k14(32'b00111110011011110011100111100011),
      .k15(32'b10111101101010101111010010011000),
      .k16(32'b00111110101011000010110110111000),
      .k17(32'b10111101110010111000000101100001),
      .k18(32'b00111101111101001010101100100110),
      .k19(32'b10111101111011111110101100011101),
      .k20(32'b00111110100000000110101010000010),
      .k21(32'b10111110100101101110001001101010),
      .k22(32'b10111110100011000100110101011101),
      .k23(32'b00111110011110110011000010011110),
      .k24(32'b00111110001010001101000001000110),
      .k25(32'b00111110100111101001100011010011),
      .k26(32'b00111110001011001110010101111010),
      .k27(32'b10111110000110000010001110010101),
      .k28(32'b10111110010010100000111110101110),
      .k29(32'b00111101010100011111101101110110),
      .k30(32'b00111110010110110010110011111001),
      .k31(32'b10111110011000111011001110100011),
      .k32(32'b10111101100101001010001111000010),
      .bias(32'b10111100000100000101011111110010)
  ) FC3 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*3-1:DATA_WIDTH*2])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110100010010100110010011111),
      .k2(32'b10111110001010011001101100011110),
      .k3(32'b00111110010010110010001110000110),
      .k4(32'b00111110010101111010100110111110),
      .k5(32'b00111101101010000110010100110100),
      .k6(32'b10111110101001111001000000011101),
      .k7(32'b00111110010111100100011101100110),
      .k8(32'b10111110100010000101001110111011),
      .k9(32'b00111110000000001000010100011010),
      .k10(32'b10111110100100010000110000100101),
      .k11(32'b00111110011101100010010001000110),
      .k12(32'b10111110001100000111001100111000),
      .k13(32'b00111101110111001111100110010000),
      .k14(32'b00111101110000011100100100000100),
      .k15(32'b10111101111100010101001111010100),
      .k16(32'b00111110101010110111010000011101),
      .k17(32'b10111101000001111000000010001000),
      .k18(32'b10111110001000000111011111111101),
      .k19(32'b10111110001110000010001111110000),
      .k20(32'b10111110100011001000011101001011),
      .k21(32'b00111101110011000110000100111000),
      .k22(32'b10111101100000001011111010110000),
      .k23(32'b10111110010010000000000011011111),
      .k24(32'b10111110011000110011110100110110),
      .k25(32'b10111110000100000100110100100011),
      .k26(32'b00111110001011101001101001000010),
      .k27(32'b00111110001011010000011001101110),
      .k28(32'b00111100010011111110000111100000),
      .k29(32'b00111110000000011011010111101010),
      .k30(32'b10111110011001011011111000001100),
      .k31(32'b00111101111100111010101111101000),
      .k32(32'b10111110100100101100000100000100),
      .bias(32'b00000000000000000000000000000000)
  ) FC4 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*4-1:DATA_WIDTH*3])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110101001011011110000100010),
      .k2(32'b00111110001100010100101100000010),
      .k3(32'b10111101110100010011111110101000),
      .k4(32'b00111110000001001010010111001010),
      .k5(32'b10111110000110101110111001001010),
      .k6(32'b10111100111110001110000110000111),
      .k7(32'b00111110010010100101011100101100),
      .k8(32'b00111110001100110100000001011100),
      .k9(32'b10111101101001111000101110010000),
      .k10(32'b10111101010110101010110011101100),
      .k11(32'b10111110000000100100100000010001),
      .k12(32'b00111110100011111110101110011011),
      .k13(32'b10111110000111111111111011000101),
      .k14(32'b00111110011011101100011110100110),
      .k15(32'b00111110100001010000010110111011),
      .k16(32'b10111101110010110001101101000111),
      .k17(32'b10111101111110110010000100101010),
      .k18(32'b00111110101001011101011010010000),
      .k19(32'b10111110001110110000101111101001),
      .k20(32'b00111110100111101111101001000101),
      .k21(32'b10111101001110111111101110110111),
      .k22(32'b10111110000100101100000001010110),
      .k23(32'b10111110101000011000000000111011),
      .k24(32'b10111110001001100100010011010110),
      .k25(32'b10111110100011011001010100000101),
      .k26(32'b10111101010111011100111010101011),
      .k27(32'b10111110011101001111110101010100),
      .k28(32'b00111110100101110010000010000111),
      .k29(32'b10111110011001111001100011010000),
      .k30(32'b00111101001000010011101110100101),
      .k31(32'b00111110011000110100110101010110),
      .k32(32'b10111110011111000111010010001011),
      .bias(32'b10111011101100100100111110110101)
  ) FC5 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*5-1:DATA_WIDTH*4])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110100101111111000111000111),
      .k2(32'b00111110101000001111100111000110),
      .k3(32'b10111110100101000000000010101101),
      .k4(32'b10111101010101010111000001110000),
      .k5(32'b00111101110001000110110000001001),
      .k6(32'b10111100000001011100110100111111),
      .k7(32'b00111110100111010100110010101010),
      .k8(32'b00111110000000100011001000110011),
      .k9(32'b10111101010010101111001110111001),
      .k10(32'b00111101110111000001100111111110),
      .k11(32'b10111110001010010011111001000000),
      .k12(32'b00111101100011101011010000110010),
      .k13(32'b10111110100000100000100110010101),
      .k14(32'b00111101011111100000101001111110),
      .k15(32'b00111101010110101001000111011111),
      .k16(32'b00111110100010001010110111111001),
      .k17(32'b10111110101101010111110000110100),
      .k18(32'b10111110010111101001101101111110),
      .k19(32'b00111110001001000111101000110111),
      .k20(32'b00111110010010100101001011010001),
      .k21(32'b10111110101011010001111001100011),
      .k22(32'b00111010110101111111010010100110),
      .k23(32'b10111101010101100111101101111010),
      .k24(32'b10111110100001101001000100001011),
      .k25(32'b10111110000000001100011011101000),
      .k26(32'b10111110001101010100010110000001),
      .k27(32'b00111110000010011000000001011111),
      .k28(32'b10111100100001011011111101110101),
      .k29(32'b10111110100100000101110110101001),
      .k30(32'b10111101111111010010000011011110),
      .k31(32'b10111110000001111111000011101100),
      .k32(32'b10111101001101000011111001101010),
      .bias(32'b10111011100110100000001010101010)
  ) FC6 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*6-1:DATA_WIDTH*5])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110100101000110010001101011),
      .k2(32'b00111110011101100110010011101010),
      .k3(32'b00111101011001001010111101110011),
      .k4(32'b00111100001101110011111100101100),
      .k5(32'b00111110100000000000101100001001),
      .k6(32'b00111110101000110000000101101001),
      .k7(32'b10111110001100011110101101011010),
      .k8(32'b10111101100000110000001101001001),
      .k9(32'b00111110001011100111011011100011),
      .k10(32'b00111110011000101111100010110100),
      .k11(32'b00111101001001110111110010010110),
      .k12(32'b00111110011000011101001100111001),
      .k13(32'b10111110010101101111110100001101),
      .k14(32'b00111110101100001101100011010101),
      .k15(32'b00111011111111110010110101011001),
      .k16(32'b10111110101000110100000011101110),
      .k17(32'b00111110100101011011000100110111),
      .k18(32'b00111110000001101101110100110110),
      .k19(32'b10111110101000000100100101100010),
      .k20(32'b10111110100001110001110100111010),
      .k21(32'b00111100101111000001100011001101),
      .k22(32'b10111110001001011010000001111010),
      .k23(32'b00111011010011010110110101010111),
      .k24(32'b00111110011110011011011011110110),
      .k25(32'b10111110100000000110000011100100),
      .k26(32'b10111110001001101110100101011101),
      .k27(32'b10111110000001001101011110010100),
      .k28(32'b10111110011101110110100100011010),
      .k29(32'b10111101010110010001001000010001),
      .k30(32'b10111110100010001010111000001100),
      .k31(32'b10111110000000001010010000111111),
      .k32(32'b10111011011110010001101011110011),
      .bias(32'b00111100010010111110011010010010)
  ) FC7 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*7-1:DATA_WIDTH*6])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111100100100001100111001001110),
      .k2(32'b10111110000001101111001101110000),
      .k3(32'b10111101010011100001110110000111),
      .k4(32'b00111110000000110000000111110011),
      .k5(32'b10111101000101100011101010000111),
      .k6(32'b00111110100001101101000001010110),
      .k7(32'b10111101111011000111001100000110),
      .k8(32'b00111100000000110011100110001101),
      .k9(32'b00111110000110100001110100010001),
      .k10(32'b00111101000010001101111000110001),
      .k11(32'b00111100100110010010011001111000),
      .k12(32'b00111110011101010001110010001111),
      .k13(32'b00111101011010011011101010110100),
      .k14(32'b00111110001110110011010011000110),
      .k15(32'b10111011011000001111000010100011),
      .k16(32'b10111110000111100011011010011111),
      .k17(32'b10111110010010111111101001011001),
      .k18(32'b10111110000001010000001000001011),
      .k19(32'b10111110000011111100101100101010),
      .k20(32'b00111101111010111011011110100011),
      .k21(32'b00111100100000011010010110010101),
      .k22(32'b00111110000001101001101110100100),
      .k23(32'b10111101010101000110110010111000),
      .k24(32'b00111101010001101000011110010101),
      .k25(32'b00111101100100100010111101100111),
      .k26(32'b00111110000000011010011111010101),
      .k27(32'b00111110011010101001010000101011),
      .k28(32'b10111110101101010001101001000011),
      .k29(32'b10111110100110010010010110110010),
      .k30(32'b10111110101101100011011101000001),
      .k31(32'b10111110100001110000010010100111),
      .k32(32'b10111110011001011011111111111010),
      .bias(32'b00111100110110000100001111000101)
  ) FC8 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*8-1:DATA_WIDTH*7])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110100001010110001001111001),
      .k2(32'b00111101111101011001110101001100),
      .k3(32'b10111101111010110010010111111100),
      .k4(32'b10111110011101011111000001011000),
      .k5(32'b10111110100011001011111011101010),
      .k6(32'b00111100101100101011110010000000),
      .k7(32'b10111110100111001011000000100101),
      .k8(32'b10111110101000101010111011111101),
      .k9(32'b10111110100010111010110111010000),
      .k10(32'b00111110100110001010011000001001),
      .k11(32'b00111110101001011001011110010001),
      .k12(32'b10111101111011110011000010110100),
      .k13(32'b10111110101000000010111001100111),
      .k14(32'b00111101111001100100111110001000),
      .k15(32'b10111101001101100011000111000000),
      .k16(32'b10111110010011110010101010011001),
      .k17(32'b00111110010110100101101101110010),
      .k18(32'b00111100111001111111101010010000),
      .k19(32'b10111100000001100111111011000000),
      .k20(32'b00111110101100010101010101100101),
      .k21(32'b10111110100010000000010110110010),
      .k22(32'b00111110100011101000001100111011),
      .k23(32'b00111110101100100111000100000101),
      .k24(32'b10111101001100111010101111111000),
      .k25(32'b00111110100010101110011100110111),
      .k26(32'b10111100100001100011110011100000),
      .k27(32'b10111110101010110111011010000111),
      .k28(32'b10111110010011010101101110000011),
      .k29(32'b10111101100011111001100011000000),
      .k30(32'b10111110100100100011110111110101),
      .k31(32'b10111110101100101011010000100111),
      .k32(32'b10111110001001000010000001101011),
      .bias(32'b00000000000000000000000000000000)
  ) FC9 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*9-1:DATA_WIDTH*8])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111101110111111010110011110011),
      .k2(32'b10111110010001101000011010110110),
      .k3(32'b10111101011101010100101001100111),
      .k4(32'b00111101101111100110110110100010),
      .k5(32'b00111100011000001101111010101110),
      .k6(32'b10111101110110100010001001000110),
      .k7(32'b00111110100011100110100001110111),
      .k8(32'b10111110100100011001110100000000),
      .k9(32'b00111110100101101011111010001000),
      .k10(32'b00111100100110110101110010010011),
      .k11(32'b10111110001100001000001000011101),
      .k12(32'b10111101100101010011111000111110),
      .k13(32'b00111110010010010110101000010111),
      .k14(32'b00111110000110010001101101000111),
      .k15(32'b00111110100110100011001100111011),
      .k16(32'b00111101101110001010001001000110),
      .k17(32'b10111110100010100101011100000000),
      .k18(32'b10111100001010011000000000100011),
      .k19(32'b10111110001100010000001010100010),
      .k20(32'b00111101111101100111100001100101),
      .k21(32'b00111110001001100111110100000110),
      .k22(32'b00111110101011011001011001110000),
      .k23(32'b10111101001000101001111110110111),
      .k24(32'b00111110101100010100111010001001),
      .k25(32'b10111110101101000111100110101111),
      .k26(32'b00111100110111110001100111100000),
      .k27(32'b00111101010001101010100001110000),
      .k28(32'b10111110011001000101110011101001),
      .k29(32'b00111110101001001111100101101111),
      .k30(32'b00111101101110111100110010001000),
      .k31(32'b00111110001111000000110101111001),
      .k32(32'b00111110100100101000010111100100),
      .bias(32'b00111100001000011001011001101000)
  ) FC10 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*10-1:DATA_WIDTH*9])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110011010010000010111111110),
      .k2(32'b00111110100001100110001001110100),
      .k3(32'b00111110100110100011100101011100),
      .k4(32'b00111110011101011000010101001001),
      .k5(32'b10111110100100010011000111111101),
      .k6(32'b00111101011100111111011011101110),
      .k7(32'b00111101011100011100011010101101),
      .k8(32'b10111110100110100110010110101101),
      .k9(32'b00111110100100001101001111110001),
      .k10(32'b00111110101001011010011001011011),
      .k11(32'b10111110000011000110010101001101),
      .k12(32'b00111110100110001000100110111110),
      .k13(32'b00111110000001101001010000011001),
      .k14(32'b00111101000111000001110001010000),
      .k15(32'b00111101000110110001001101110001),
      .k16(32'b00111101100110110101011001110111),
      .k17(32'b00111110100110010100101000101101),
      .k18(32'b10111110010111001111100001001011),
      .k19(32'b10111101001111100011100110001010),
      .k20(32'b00111110000000011111100010011000),
      .k21(32'b00111110001001011011100000011111),
      .k22(32'b10111110011110101110110110100100),
      .k23(32'b10111110001110100010010001110100),
      .k24(32'b00111110001111101010111110110110),
      .k25(32'b10111101001101110110010000011010),
      .k26(32'b10111101111000010110000000111110),
      .k27(32'b10111101001101111111111110010000),
      .k28(32'b10111110000110011010101000010010),
      .k29(32'b00111110011000010010010100001100),
      .k30(32'b00111110001100110110100000110011),
      .k31(32'b10111110010001110010111001100110),
      .k32(32'b00111101010111100011000100010001),
      .bias(32'b00111100001001110011000111110000)
  ) FC11 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*11-1:DATA_WIDTH*10])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110001001110100000011001010),
      .k2(32'b00111110101011000010011100000001),
      .k3(32'b00111110101000011111000111101100),
      .k4(32'b10111110000000001010011001001010),
      .k5(32'b00111110100100110010001010000011),
      .k6(32'b00111110101100010101101001100001),
      .k7(32'b00111110011011010001001011111001),
      .k8(32'b00111110001110000001100101101101),
      .k9(32'b10111110000010101011110010100110),
      .k10(32'b00111100101100011111000111100000),
      .k11(32'b00111100110100010001100111100110),
      .k12(32'b10111110010110101101101010110000),
      .k13(32'b10111101001100000010110101110101),
      .k14(32'b00111110000100100101110011001110),
      .k15(32'b00111101111111001100110011100010),
      .k16(32'b00111110100100110110011000001011),
      .k17(32'b10111110010011010111010110010100),
      .k18(32'b00111110001011100000100100111010),
      .k19(32'b00111101010100010100001110110001),
      .k20(32'b00111101001000001011000010011000),
      .k21(32'b00111110101010011111000100000011),
      .k22(32'b00111100100000000111001010001101),
      .k23(32'b10111110100011011111010111001110),
      .k24(32'b10111110100001000101111010010100),
      .k25(32'b10111110101100011111111011010001),
      .k26(32'b00111110101011110111001011100000),
      .k27(32'b10111101100101110111100001000100),
      .k28(32'b00111110001101100011001011001100),
      .k29(32'b00111110010011010100000110101101),
      .k30(32'b10111110000011001111101101101101),
      .k31(32'b10111110101011001011110000000111),
      .k32(32'b10111110100011111011111101111000),
      .bias(32'b10111100000110001000100011110000)
  ) FC12 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*12-1:DATA_WIDTH*11])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110100011000011000000110001),
      .k2(32'b10111101100010000010101101011000),
      .k3(32'b00111110011000001101010110011010),
      .k4(32'b10111110000100000010000011010101),
      .k5(32'b10111110000110111011001101101111),
      .k6(32'b00111101001011110000110111100000),
      .k7(32'b10111110000100100110010000010110),
      .k8(32'b10111110011000000010011111110010),
      .k9(32'b00111100010000001101010110100000),
      .k10(32'b10111110101001111010111010010110),
      .k11(32'b10111110011100101111000011110000),
      .k12(32'b00111110000101110110111110010010),
      .k13(32'b10111101101010101111101110011000),
      .k14(32'b10111101111010000111100110001110),
      .k15(32'b10111110100001101100101011111010),
      .k16(32'b10111110011001100001101101101000),
      .k17(32'b10111110100010010110001101001011),
      .k18(32'b10111110100110101010101111010000),
      .k19(32'b00111110100010011110010110000101),
      .k20(32'b10111101000010001010011111011000),
      .k21(32'b10111101110001001010011110011100),
      .k22(32'b00111110011100010101001110010110),
      .k23(32'b00111110101001011101111000010011),
      .k24(32'b00111101110101100111100000110000),
      .k25(32'b10111110000010011011000110110111),
      .k26(32'b00111110101010011000111100010001),
      .k27(32'b00111110011001100110011011011110),
      .k28(32'b10111101100011101010111010010100),
      .k29(32'b00111110010110100001000011010010),
      .k30(32'b10111110011110100111010111100110),
      .k31(32'b00111100110000110000101111010000),
      .k32(32'b10111110010110011010000011110001),
      .bias(32'b00000000000000000000000000000000)
  ) FC13 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*13-1:DATA_WIDTH*12])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111100101011010101010011011101),
      .k2(32'b10111110101000110111101101010110),
      .k3(32'b00111101101000000001101111100100),
      .k4(32'b10111110011000000010111110111001),
      .k5(32'b10111110010100110011111010110101),
      .k6(32'b10111110000001111001110011010000),
      .k7(32'b00111110010110110111111111101101),
      .k8(32'b00111110000000000011101100110010),
      .k9(32'b00111101001110000101000101001011),
      .k10(32'b00111110101101010100100100111001),
      .k11(32'b10111110001100010010101110000000),
      .k12(32'b10111110100000011011101101111101),
      .k13(32'b10111110100101100010111111010111),
      .k14(32'b00111110001101001000010000000100),
      .k15(32'b10111110000110111101010011010000),
      .k16(32'b00111011111100011101001001011001),
      .k17(32'b00111110101011001011110100010101),
      .k18(32'b00111101101100111100110011101001),
      .k19(32'b00111101110010011000101101011010),
      .k20(32'b00111110101010010110100011101011),
      .k21(32'b00111110001001101100111000110000),
      .k22(32'b00111110101001101110000101110001),
      .k23(32'b10111100011101011010100100111011),
      .k24(32'b10111110101010101101110111001011),
      .k25(32'b10111110000111011101001110101110),
      .k26(32'b10111110010010011001000110001101),
      .k27(32'b10111101100011011011111000101100),
      .k28(32'b00111110011100101111001111011110),
      .k29(32'b10111110100010001000010011001100),
      .k30(32'b00111110101011101110100010000001),
      .k31(32'b10111110011011001100011011100001),
      .k32(32'b10111110100011010011110100111000),
      .bias(32'b00111011001101111100010000010100)
  ) FC14 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*14-1:DATA_WIDTH*13])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b10111110100111111110011110110000),
      .k2(32'b00111101100111001111011001011001),
      .k3(32'b10111110100011110000011000011011),
      .k4(32'b00111110101100001111110100010100),
      .k5(32'b10111110011100001000111110101010),
      .k6(32'b00111100101101101100000100010010),
      .k7(32'b10111110100010011001000111101010),
      .k8(32'b00111110100101110100111111101010),
      .k9(32'b00111110010001100010001011100111),
      .k10(32'b10111101111011011011011100011011),
      .k11(32'b10111110101010001010100111011010),
      .k12(32'b10111110100101100000000110101111),
      .k13(32'b10111101110010110000011001101101),
      .k14(32'b10111110010001010110100011101010),
      .k15(32'b00111101000110000101101110101101),
      .k16(32'b10111110001000000110100010000011),
      .k17(32'b00111110000111000011110011001000),
      .k18(32'b00111110100100100010001011001111),
      .k19(32'b00111101100100001011000001010011),
      .k20(32'b10111101111000001011010111011100),
      .k21(32'b00111110000000000000000000001010),
      .k22(32'b10111110100001110100000011010101),
      .k23(32'b00111110100111010011010001100001),
      .k24(32'b00111101100001010001111111110010),
      .k25(32'b00111101010001110101000100000001),
      .k26(32'b00111110100111101010101011100010),
      .k27(32'b10111110001001011100001010110000),
      .k28(32'b00111110100101100100000101010110),
      .k29(32'b00111101001101101100101100110111),
      .k30(32'b10111110011001001010011011011100),
      .k31(32'b00111110011010001001100000101011),
      .k32(32'b00111110100010110001111000000111),
      .bias(32'b00111100010101011111011000100100)
  ) FC15 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*15-1:DATA_WIDTH*14])  
  );

  FC#(
      .DATA_WIDTH(DATA_WIDTH),
      .k1(32'b00111110000101110001100000110010),
      .k2(32'b00111100111001101001010011110000),
      .k3(32'b10111110000110011111001101110101),
      .k4(32'b10111101110100111001011100100000),
      .k5(32'b10111101110111010100001000101100),
      .k6(32'b10111101101111010011000101110100),
      .k7(32'b10111110100011110100000001010110),
      .k8(32'b00111110101010110011001110110101),
      .k9(32'b00111101101110110000100001110100),
      .k10(32'b00111011111101001101000111000000),
      .k11(32'b00111110000100010011011001101010),
      .k12(32'b10111110100110000101010010001000),
      .k13(32'b00111101101100111001000101101000),
      .k14(32'b10111110101001001001100100000011),
      .k15(32'b10111110101100111110001101100110),
      .k16(32'b10111110000000001100001110001101),
      .k17(32'b00111101101010101100010100111100),
      .k18(32'b10111101011110000100100111010000),
      .k19(32'b10111110100100101001000001110100),
      .k20(32'b10111110010001010011011101010000),
      .k21(32'b00111110000110101101110000001110),
      .k22(32'b00111110101001011000010101011101),
      .k23(32'b10111110100001001000100110111100),
      .k24(32'b10111110010001011100100101100110),
      .k25(32'b10111110100101101100011101111010),
      .k26(32'b00111110001101110010000101000110),
      .k27(32'b10111110100010010011100111010100),
      .k28(32'b00111110001100011011101111100010),
      .k29(32'b00111100001000011100101110000000),
      .k30(32'b10111110010101111010011111100100),
      .k31(32'b10111110101011010100110010111110),
      .k32(32'b00111110101010000110111010101101),
      .bias(32'b00000000000000000000000000000000)
  ) FC16 (
      .i_data(i_data[DATA_WIDTH*32-1:0]),
      .clk(clk), 
      .rst(rst), 
      .valid_in(valid_in),
      .valid_pipeline_FC(valid_pipeline_FC),
      .o_data(o_data[DATA_WIDTH*16-1:DATA_WIDTH*15])  
  );

 control_FC control(
       .valid_in_FC(valid_in), 
       .clk(clk), 
       .rst(rst),
       .valid_out(valid_out),
       .valid_in_FC1(valid_pipeline_FC)  
  );
endmodule
